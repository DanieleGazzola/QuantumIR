module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644;
  assign n65 = x0 & x32;
  assign n67 = ~x32 & x33;
  assign n68 = ~x0 & n67;
  assign n70 = x32 & ~x33;
  assign n69 = x32 & x33;
  assign n71 = n70 ^ n69;
  assign n72 = n69 ^ x1;
  assign n73 = n72 ^ n69;
  assign n74 = n71 & n73;
  assign n75 = n74 ^ n69;
  assign n76 = ~n68 & ~n75;
  assign n66 = x33 & ~n65;
  assign n77 = n76 ^ n66;
  assign n81 = ~x1 & n67;
  assign n82 = n69 ^ x2;
  assign n83 = n82 ^ n69;
  assign n84 = n71 & n83;
  assign n85 = n84 ^ n69;
  assign n86 = ~n81 & ~n85;
  assign n79 = x34 ^ x33;
  assign n80 = x0 & n79;
  assign n87 = n86 ^ n80;
  assign n78 = n66 & ~n76;
  assign n88 = n87 ^ n78;
  assign n114 = n80 ^ n78;
  assign n115 = n87 & n114;
  assign n116 = n115 ^ n78;
  assign n106 = ~x2 & n67;
  assign n107 = n69 ^ x3;
  assign n108 = n107 ^ n69;
  assign n109 = n71 & n108;
  assign n110 = n109 ^ n69;
  assign n111 = ~n106 & ~n110;
  assign n102 = x33 ^ x0;
  assign n103 = ~n79 & n102;
  assign n104 = n103 ^ x0;
  assign n105 = x35 & ~n104;
  assign n112 = n111 ^ n105;
  assign n89 = x35 & n79;
  assign n90 = ~x1 & n89;
  assign n91 = x35 ^ x34;
  assign n92 = ~n79 & n91;
  assign n93 = x35 & n92;
  assign n94 = ~x0 & n93;
  assign n95 = ~n90 & ~n94;
  assign n96 = ~x35 & n79;
  assign n97 = x1 & n96;
  assign n98 = ~x35 & n92;
  assign n99 = x0 & n98;
  assign n100 = ~n97 & ~n99;
  assign n101 = n95 & n100;
  assign n113 = n112 ^ n101;
  assign n117 = n116 ^ n113;
  assign n137 = n116 ^ n101;
  assign n138 = ~n113 & ~n137;
  assign n139 = n138 ^ n116;
  assign n129 = ~x3 & n67;
  assign n130 = n69 ^ x4;
  assign n131 = n130 ^ n69;
  assign n132 = n71 & n131;
  assign n133 = n132 ^ n69;
  assign n134 = ~n129 & ~n133;
  assign n121 = x2 & n96;
  assign n122 = x1 & n98;
  assign n123 = ~n121 & ~n122;
  assign n124 = ~x2 & n89;
  assign n125 = ~x1 & n93;
  assign n126 = ~n124 & ~n125;
  assign n127 = n123 & n126;
  assign n119 = x36 ^ x35;
  assign n120 = x0 & n119;
  assign n128 = n127 ^ n120;
  assign n135 = n134 ^ n128;
  assign n118 = n105 & ~n111;
  assign n136 = n135 ^ n118;
  assign n140 = n139 ^ n136;
  assign n179 = n139 ^ n118;
  assign n180 = ~n136 & n179;
  assign n181 = n180 ^ n139;
  assign n174 = n134 ^ n120;
  assign n175 = n134 ^ n127;
  assign n176 = ~n174 & ~n175;
  assign n177 = n176 ^ n120;
  assign n159 = x37 & n119;
  assign n160 = ~x1 & n159;
  assign n161 = x37 ^ x36;
  assign n162 = ~n119 & n161;
  assign n163 = x37 & n162;
  assign n164 = ~x0 & n163;
  assign n165 = ~n160 & ~n164;
  assign n166 = ~x37 & n119;
  assign n167 = x1 & n166;
  assign n168 = ~x37 & n162;
  assign n169 = x0 & n168;
  assign n170 = ~n167 & ~n169;
  assign n171 = n165 & n170;
  assign n152 = x3 & n96;
  assign n153 = x2 & n98;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~x3 & n89;
  assign n156 = ~x2 & n93;
  assign n157 = ~n155 & ~n156;
  assign n158 = n154 & n157;
  assign n172 = n171 ^ n158;
  assign n145 = ~x4 & n67;
  assign n146 = n69 ^ x5;
  assign n147 = n146 ^ n69;
  assign n148 = n71 & n147;
  assign n149 = n148 ^ n69;
  assign n150 = ~n145 & ~n149;
  assign n141 = x35 ^ x0;
  assign n142 = ~n119 & n141;
  assign n143 = n142 ^ x0;
  assign n144 = x37 & ~n143;
  assign n151 = n150 ^ n144;
  assign n173 = n172 ^ n151;
  assign n178 = n177 ^ n173;
  assign n182 = n181 ^ n178;
  assign n214 = n181 ^ n173;
  assign n215 = n178 & ~n214;
  assign n216 = n215 ^ n181;
  assign n210 = n171 ^ n151;
  assign n211 = n172 & ~n210;
  assign n212 = n211 ^ n158;
  assign n207 = n144 & ~n150;
  assign n200 = ~x2 & n159;
  assign n201 = ~x1 & n163;
  assign n202 = ~n200 & ~n201;
  assign n203 = x2 & n166;
  assign n204 = x1 & n168;
  assign n205 = ~n203 & ~n204;
  assign n206 = n202 & n205;
  assign n208 = n207 ^ n206;
  assign n192 = ~x4 & n89;
  assign n193 = ~x3 & n93;
  assign n194 = ~n192 & ~n193;
  assign n195 = x4 & n96;
  assign n196 = x3 & n98;
  assign n197 = ~n195 & ~n196;
  assign n198 = n194 & n197;
  assign n185 = ~x5 & n67;
  assign n186 = n69 ^ x6;
  assign n187 = n186 ^ n69;
  assign n188 = n71 & n187;
  assign n189 = n188 ^ n69;
  assign n190 = ~n185 & ~n189;
  assign n183 = x38 ^ x37;
  assign n184 = x0 & n183;
  assign n191 = n190 ^ n184;
  assign n199 = n198 ^ n191;
  assign n209 = n208 ^ n199;
  assign n213 = n212 ^ n209;
  assign n217 = n216 ^ n213;
  assign n267 = n216 ^ n209;
  assign n268 = ~n213 & ~n267;
  assign n269 = n268 ^ n216;
  assign n263 = n207 ^ n199;
  assign n264 = ~n208 & ~n263;
  assign n265 = n264 ^ n206;
  assign n258 = n198 ^ n190;
  assign n259 = ~n191 & ~n258;
  assign n260 = n259 ^ n184;
  assign n251 = ~x6 & n67;
  assign n252 = n69 ^ x7;
  assign n253 = n252 ^ n69;
  assign n254 = n71 & n253;
  assign n255 = n254 ^ n69;
  assign n256 = ~n251 & ~n255;
  assign n247 = x37 ^ x0;
  assign n248 = ~n183 & n247;
  assign n249 = n248 ^ x0;
  assign n250 = x39 & ~n249;
  assign n257 = n256 ^ n250;
  assign n261 = n260 ^ n257;
  assign n238 = x5 & n96;
  assign n239 = x4 & n98;
  assign n240 = ~n238 & ~n239;
  assign n241 = ~x5 & n89;
  assign n242 = ~x4 & n93;
  assign n243 = ~n241 & ~n242;
  assign n244 = n240 & n243;
  assign n225 = x39 & n183;
  assign n226 = ~x1 & n225;
  assign n227 = x39 ^ x38;
  assign n228 = ~n183 & n227;
  assign n229 = x39 & n228;
  assign n230 = ~x0 & n229;
  assign n231 = ~n226 & ~n230;
  assign n232 = ~x39 & n183;
  assign n233 = x1 & n232;
  assign n234 = ~x39 & n228;
  assign n235 = x0 & n234;
  assign n236 = ~n233 & ~n235;
  assign n237 = n231 & n236;
  assign n245 = n244 ^ n237;
  assign n218 = x3 & n166;
  assign n219 = x2 & n168;
  assign n220 = ~n218 & ~n219;
  assign n221 = ~x3 & n159;
  assign n222 = ~x2 & n163;
  assign n223 = ~n221 & ~n222;
  assign n224 = n220 & n223;
  assign n246 = n245 ^ n224;
  assign n262 = n261 ^ n246;
  assign n266 = n265 ^ n262;
  assign n270 = n269 ^ n266;
  assign n316 = n269 ^ n262;
  assign n317 = n266 & n316;
  assign n318 = n317 ^ n269;
  assign n311 = n257 ^ n246;
  assign n312 = n260 ^ n246;
  assign n313 = n311 & n312;
  assign n314 = n313 ^ n257;
  assign n305 = n237 ^ n224;
  assign n306 = n244 ^ n224;
  assign n307 = n305 & ~n306;
  assign n308 = n307 ^ n237;
  assign n297 = ~x2 & n225;
  assign n298 = ~x1 & n229;
  assign n299 = ~n297 & ~n298;
  assign n300 = x2 & n232;
  assign n301 = x1 & n234;
  assign n302 = ~n300 & ~n301;
  assign n303 = n299 & n302;
  assign n290 = ~x7 & n67;
  assign n291 = n69 ^ x8;
  assign n292 = n291 ^ n69;
  assign n293 = n71 & n292;
  assign n294 = n293 ^ n69;
  assign n295 = ~n290 & ~n294;
  assign n288 = x40 ^ x39;
  assign n289 = x0 & n288;
  assign n296 = n295 ^ n289;
  assign n304 = n303 ^ n296;
  assign n309 = n308 ^ n304;
  assign n279 = ~x4 & n159;
  assign n280 = ~x3 & n163;
  assign n281 = ~n279 & ~n280;
  assign n282 = x4 & n166;
  assign n283 = x3 & n168;
  assign n284 = ~n282 & ~n283;
  assign n285 = n281 & n284;
  assign n272 = ~x6 & n89;
  assign n273 = ~x5 & n93;
  assign n274 = ~n272 & ~n273;
  assign n275 = x6 & n96;
  assign n276 = x5 & n98;
  assign n277 = ~n275 & ~n276;
  assign n278 = n274 & n277;
  assign n286 = n285 ^ n278;
  assign n271 = n250 & ~n256;
  assign n287 = n286 ^ n271;
  assign n310 = n309 ^ n287;
  assign n315 = n314 ^ n310;
  assign n319 = n318 ^ n315;
  assign n382 = n318 ^ n310;
  assign n383 = ~n315 & ~n382;
  assign n384 = n383 ^ n318;
  assign n377 = n304 ^ n287;
  assign n378 = n308 ^ n287;
  assign n379 = n377 & n378;
  assign n380 = n379 ^ n304;
  assign n372 = n285 ^ n271;
  assign n373 = n286 & n372;
  assign n374 = n373 ^ n278;
  assign n365 = ~x8 & n67;
  assign n366 = n69 ^ x9;
  assign n367 = n366 ^ n69;
  assign n368 = n71 & n367;
  assign n369 = n368 ^ n69;
  assign n370 = ~n365 & ~n369;
  assign n357 = ~x3 & n225;
  assign n358 = ~x2 & n229;
  assign n359 = ~n357 & ~n358;
  assign n360 = x3 & n232;
  assign n361 = x2 & n234;
  assign n362 = ~n360 & ~n361;
  assign n363 = n359 & n362;
  assign n344 = x41 & n288;
  assign n345 = ~x1 & n344;
  assign n346 = x41 ^ x40;
  assign n347 = ~n288 & n346;
  assign n348 = x41 & n347;
  assign n349 = ~x0 & n348;
  assign n350 = ~n345 & ~n349;
  assign n351 = ~x41 & n288;
  assign n352 = x1 & n351;
  assign n353 = ~x41 & n347;
  assign n354 = x0 & n353;
  assign n355 = ~n352 & ~n354;
  assign n356 = n350 & n355;
  assign n364 = n363 ^ n356;
  assign n371 = n370 ^ n364;
  assign n375 = n374 ^ n371;
  assign n340 = n303 ^ n295;
  assign n341 = ~n296 & ~n340;
  assign n342 = n341 ^ n289;
  assign n331 = ~x7 & n89;
  assign n332 = ~x6 & n93;
  assign n333 = ~n331 & ~n332;
  assign n334 = x7 & n96;
  assign n335 = x6 & n98;
  assign n336 = ~n334 & ~n335;
  assign n337 = n333 & n336;
  assign n327 = x39 ^ x0;
  assign n328 = ~n288 & n327;
  assign n329 = n328 ^ x0;
  assign n330 = x41 & ~n329;
  assign n338 = n337 ^ n330;
  assign n320 = x5 & n166;
  assign n321 = x4 & n168;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~x5 & n159;
  assign n324 = ~x4 & n163;
  assign n325 = ~n323 & ~n324;
  assign n326 = n322 & n325;
  assign n339 = n338 ^ n326;
  assign n343 = n342 ^ n339;
  assign n376 = n375 ^ n343;
  assign n381 = n380 ^ n376;
  assign n385 = n384 ^ n381;
  assign n442 = n384 ^ n376;
  assign n443 = ~n381 & n442;
  assign n444 = n443 ^ n384;
  assign n437 = n371 ^ n343;
  assign n438 = n374 ^ n343;
  assign n439 = ~n437 & n438;
  assign n440 = n439 ^ n371;
  assign n432 = n342 ^ n338;
  assign n433 = n339 & n432;
  assign n434 = n433 ^ n326;
  assign n424 = ~x9 & n67;
  assign n425 = n69 ^ x10;
  assign n426 = n425 ^ n69;
  assign n427 = n71 & n426;
  assign n428 = n427 ^ n69;
  assign n429 = ~n424 & ~n428;
  assign n417 = ~x2 & n344;
  assign n418 = ~x1 & n348;
  assign n419 = ~n417 & ~n418;
  assign n420 = x2 & n351;
  assign n421 = x1 & n353;
  assign n422 = ~n420 & ~n421;
  assign n423 = n419 & n422;
  assign n430 = n429 ^ n423;
  assign n410 = ~x6 & n159;
  assign n411 = ~x5 & n163;
  assign n412 = ~n410 & ~n411;
  assign n413 = x6 & n166;
  assign n414 = x5 & n168;
  assign n415 = ~n413 & ~n414;
  assign n416 = n412 & n415;
  assign n431 = n430 ^ n416;
  assign n435 = n434 ^ n431;
  assign n405 = n370 ^ n356;
  assign n406 = ~n364 & n405;
  assign n407 = n406 ^ n370;
  assign n404 = n330 & ~n337;
  assign n408 = n407 ^ n404;
  assign n395 = ~x8 & n89;
  assign n396 = ~x7 & n93;
  assign n397 = ~n395 & ~n396;
  assign n398 = x8 & n96;
  assign n399 = x7 & n98;
  assign n400 = ~n398 & ~n399;
  assign n401 = n397 & n400;
  assign n393 = x42 ^ x41;
  assign n394 = x0 & n393;
  assign n402 = n401 ^ n394;
  assign n386 = x4 & n232;
  assign n387 = x3 & n234;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~x4 & n225;
  assign n390 = ~x3 & n229;
  assign n391 = ~n389 & ~n390;
  assign n392 = n388 & n391;
  assign n403 = n402 ^ n392;
  assign n409 = n408 ^ n403;
  assign n436 = n435 ^ n409;
  assign n441 = n440 ^ n436;
  assign n445 = n444 ^ n441;
  assign n520 = n444 ^ n436;
  assign n521 = ~n441 & ~n520;
  assign n522 = n521 ^ n444;
  assign n515 = n431 ^ n409;
  assign n516 = n434 ^ n409;
  assign n517 = n515 & ~n516;
  assign n518 = n517 ^ n431;
  assign n511 = n404 ^ n403;
  assign n512 = n408 & n511;
  assign n513 = n512 ^ n403;
  assign n502 = ~x10 & n67;
  assign n503 = n69 ^ x11;
  assign n504 = n503 ^ n69;
  assign n505 = n71 & n504;
  assign n506 = n505 ^ n69;
  assign n507 = ~n502 & ~n506;
  assign n494 = ~x3 & n344;
  assign n495 = ~x2 & n348;
  assign n496 = ~n494 & ~n495;
  assign n497 = x3 & n351;
  assign n498 = x2 & n353;
  assign n499 = ~n497 & ~n498;
  assign n500 = n496 & n499;
  assign n487 = ~x5 & n225;
  assign n488 = ~x4 & n229;
  assign n489 = ~n487 & ~n488;
  assign n490 = x5 & n232;
  assign n491 = x4 & n234;
  assign n492 = ~n490 & ~n491;
  assign n493 = n489 & n492;
  assign n501 = n500 ^ n493;
  assign n508 = n507 ^ n501;
  assign n483 = n401 ^ n392;
  assign n484 = ~n402 & ~n483;
  assign n485 = n484 ^ n394;
  assign n480 = n423 ^ n416;
  assign n481 = n430 & ~n480;
  assign n482 = n481 ^ n429;
  assign n486 = n485 ^ n482;
  assign n509 = n508 ^ n486;
  assign n471 = x9 & n96;
  assign n472 = x8 & n98;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~x9 & n89;
  assign n475 = ~x8 & n93;
  assign n476 = ~n474 & ~n475;
  assign n477 = n473 & n476;
  assign n467 = x41 ^ x0;
  assign n468 = ~n393 & n467;
  assign n469 = n468 ^ x0;
  assign n470 = x43 & ~n469;
  assign n478 = n477 ^ n470;
  assign n453 = ~x43 & n393;
  assign n454 = x1 & n453;
  assign n455 = x43 ^ x42;
  assign n456 = ~n393 & n455;
  assign n457 = ~x43 & n456;
  assign n458 = x0 & n457;
  assign n459 = ~n454 & ~n458;
  assign n460 = x43 & n393;
  assign n461 = ~x1 & n460;
  assign n462 = x43 & n456;
  assign n463 = ~x0 & n462;
  assign n464 = ~n461 & ~n463;
  assign n465 = n459 & n464;
  assign n446 = ~x7 & n159;
  assign n447 = ~x6 & n163;
  assign n448 = ~n446 & ~n447;
  assign n449 = x7 & n166;
  assign n450 = x6 & n168;
  assign n451 = ~n449 & ~n450;
  assign n452 = n448 & n451;
  assign n466 = n465 ^ n452;
  assign n479 = n478 ^ n466;
  assign n510 = n509 ^ n479;
  assign n514 = n513 ^ n510;
  assign n519 = n518 ^ n514;
  assign n523 = n522 ^ n519;
  assign n591 = n522 ^ n514;
  assign n592 = ~n519 & ~n591;
  assign n593 = n592 ^ n522;
  assign n587 = n513 ^ n509;
  assign n588 = ~n510 & ~n587;
  assign n589 = n588 ^ n479;
  assign n582 = n508 ^ n482;
  assign n583 = n486 & n582;
  assign n584 = n583 ^ n508;
  assign n578 = n507 ^ n493;
  assign n579 = ~n501 & n578;
  assign n580 = n579 ^ n507;
  assign n576 = n470 & ~n477;
  assign n569 = ~x8 & n159;
  assign n570 = ~x7 & n163;
  assign n571 = ~n569 & ~n570;
  assign n572 = x8 & n166;
  assign n573 = x7 & n168;
  assign n574 = ~n572 & ~n573;
  assign n575 = n571 & n574;
  assign n577 = n576 ^ n575;
  assign n581 = n580 ^ n577;
  assign n585 = n584 ^ n581;
  assign n565 = n478 ^ n465;
  assign n566 = n466 & ~n565;
  assign n567 = n566 ^ n452;
  assign n556 = ~x11 & n67;
  assign n557 = n69 ^ x12;
  assign n558 = n557 ^ n69;
  assign n559 = n71 & n558;
  assign n560 = n559 ^ n69;
  assign n561 = ~n556 & ~n560;
  assign n549 = ~x4 & n344;
  assign n550 = ~x3 & n348;
  assign n551 = ~n549 & ~n550;
  assign n552 = x4 & n351;
  assign n553 = x3 & n353;
  assign n554 = ~n552 & ~n553;
  assign n555 = n551 & n554;
  assign n562 = n561 ^ n555;
  assign n542 = x2 & n453;
  assign n543 = x1 & n457;
  assign n544 = ~n542 & ~n543;
  assign n545 = ~x2 & n460;
  assign n546 = ~x1 & n462;
  assign n547 = ~n545 & ~n546;
  assign n548 = n544 & n547;
  assign n563 = n562 ^ n548;
  assign n533 = x10 & n96;
  assign n534 = x9 & n98;
  assign n535 = ~n533 & ~n534;
  assign n536 = ~x10 & n89;
  assign n537 = ~x9 & n93;
  assign n538 = ~n536 & ~n537;
  assign n539 = n535 & n538;
  assign n531 = x44 ^ x43;
  assign n532 = x0 & n531;
  assign n540 = n539 ^ n532;
  assign n524 = ~x6 & n225;
  assign n525 = ~x5 & n229;
  assign n526 = ~n524 & ~n525;
  assign n527 = x6 & n232;
  assign n528 = x5 & n234;
  assign n529 = ~n527 & ~n528;
  assign n530 = n526 & n529;
  assign n541 = n540 ^ n530;
  assign n564 = n563 ^ n541;
  assign n568 = n567 ^ n564;
  assign n586 = n585 ^ n568;
  assign n590 = n589 ^ n586;
  assign n594 = n593 ^ n590;
  assign n681 = n593 ^ n586;
  assign n682 = ~n590 & ~n681;
  assign n683 = n682 ^ n593;
  assign n677 = n581 ^ n568;
  assign n678 = n585 & n677;
  assign n679 = n678 ^ n568;
  assign n672 = n567 ^ n563;
  assign n673 = ~n564 & ~n672;
  assign n674 = n673 ^ n541;
  assign n668 = n555 ^ n548;
  assign n669 = n562 & ~n668;
  assign n670 = n669 ^ n561;
  assign n663 = n532 ^ n530;
  assign n664 = n539 ^ n530;
  assign n665 = ~n663 & ~n664;
  assign n666 = n665 ^ n532;
  assign n656 = ~x12 & n67;
  assign n657 = n69 ^ x13;
  assign n658 = n657 ^ n69;
  assign n659 = n71 & n658;
  assign n660 = n659 ^ n69;
  assign n661 = ~n656 & ~n660;
  assign n652 = x43 ^ x0;
  assign n653 = ~n531 & n652;
  assign n654 = n653 ^ x0;
  assign n655 = x45 & ~n654;
  assign n662 = n661 ^ n655;
  assign n667 = n666 ^ n662;
  assign n671 = n670 ^ n667;
  assign n675 = n674 ^ n671;
  assign n648 = n580 ^ n576;
  assign n649 = ~n577 & n648;
  assign n650 = n649 ^ n575;
  assign n638 = x3 & n453;
  assign n639 = x2 & n457;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~x3 & n460;
  assign n642 = ~x2 & n462;
  assign n643 = ~n641 & ~n642;
  assign n644 = n640 & n643;
  assign n631 = ~x9 & n159;
  assign n632 = ~x8 & n163;
  assign n633 = ~n631 & ~n632;
  assign n634 = x9 & n166;
  assign n635 = x8 & n168;
  assign n636 = ~n634 & ~n635;
  assign n637 = n633 & n636;
  assign n645 = n644 ^ n637;
  assign n618 = x45 & n531;
  assign n619 = ~x1 & n618;
  assign n620 = x45 ^ x44;
  assign n621 = ~n531 & n620;
  assign n622 = x45 & n621;
  assign n623 = ~x0 & n622;
  assign n624 = ~n619 & ~n623;
  assign n625 = ~x45 & n531;
  assign n626 = x1 & n625;
  assign n627 = ~x45 & n621;
  assign n628 = x0 & n627;
  assign n629 = ~n626 & ~n628;
  assign n630 = n624 & n629;
  assign n646 = n645 ^ n630;
  assign n609 = ~x11 & n89;
  assign n610 = ~x10 & n93;
  assign n611 = ~n609 & ~n610;
  assign n612 = x11 & n96;
  assign n613 = x10 & n98;
  assign n614 = ~n612 & ~n613;
  assign n615 = n611 & n614;
  assign n602 = x7 & n232;
  assign n603 = x6 & n234;
  assign n604 = ~n602 & ~n603;
  assign n605 = ~x7 & n225;
  assign n606 = ~x6 & n229;
  assign n607 = ~n605 & ~n606;
  assign n608 = n604 & n607;
  assign n616 = n615 ^ n608;
  assign n595 = x5 & n351;
  assign n596 = x4 & n353;
  assign n597 = ~n595 & ~n596;
  assign n598 = ~x5 & n344;
  assign n599 = ~x4 & n348;
  assign n600 = ~n598 & ~n599;
  assign n601 = n597 & n600;
  assign n617 = n616 ^ n601;
  assign n647 = n646 ^ n617;
  assign n651 = n650 ^ n647;
  assign n676 = n675 ^ n651;
  assign n680 = n679 ^ n676;
  assign n684 = n683 ^ n680;
  assign n764 = n683 ^ n676;
  assign n765 = n680 & ~n764;
  assign n766 = n765 ^ n683;
  assign n760 = n674 ^ n651;
  assign n761 = n675 & n760;
  assign n762 = n761 ^ n671;
  assign n756 = n650 ^ n646;
  assign n757 = n647 & ~n756;
  assign n758 = n757 ^ n617;
  assign n751 = n670 ^ n666;
  assign n752 = ~n667 & n751;
  assign n753 = n752 ^ n662;
  assign n741 = x2 & n625;
  assign n742 = x1 & n627;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~x2 & n618;
  assign n745 = ~x1 & n622;
  assign n746 = ~n744 & ~n745;
  assign n747 = n743 & n746;
  assign n734 = x4 & n453;
  assign n735 = x3 & n457;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~x4 & n460;
  assign n738 = ~x3 & n462;
  assign n739 = ~n737 & ~n738;
  assign n740 = n736 & n739;
  assign n748 = n747 ^ n740;
  assign n733 = n655 & ~n661;
  assign n749 = n748 ^ n733;
  assign n724 = ~x6 & n344;
  assign n725 = ~x5 & n348;
  assign n726 = ~n724 & ~n725;
  assign n727 = x6 & n351;
  assign n728 = x5 & n353;
  assign n729 = ~n727 & ~n728;
  assign n730 = n726 & n729;
  assign n717 = x8 & n232;
  assign n718 = x7 & n234;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~x8 & n225;
  assign n721 = ~x7 & n229;
  assign n722 = ~n720 & ~n721;
  assign n723 = n719 & n722;
  assign n731 = n730 ^ n723;
  assign n710 = x10 & n166;
  assign n711 = x9 & n168;
  assign n712 = ~n710 & ~n711;
  assign n713 = ~x10 & n159;
  assign n714 = ~x9 & n163;
  assign n715 = ~n713 & ~n714;
  assign n716 = n712 & n715;
  assign n732 = n731 ^ n716;
  assign n750 = n749 ^ n732;
  assign n754 = n753 ^ n750;
  assign n705 = n644 ^ n630;
  assign n706 = n645 & ~n705;
  assign n707 = n706 ^ n637;
  assign n702 = n615 ^ n601;
  assign n703 = n616 & ~n702;
  assign n704 = n703 ^ n608;
  assign n708 = n707 ^ n704;
  assign n694 = ~x12 & n89;
  assign n695 = ~x11 & n93;
  assign n696 = ~n694 & ~n695;
  assign n697 = x12 & n96;
  assign n698 = x11 & n98;
  assign n699 = ~n697 & ~n698;
  assign n700 = n696 & n699;
  assign n687 = ~x13 & n67;
  assign n688 = n69 ^ x14;
  assign n689 = n688 ^ n69;
  assign n690 = n71 & n689;
  assign n691 = n690 ^ n69;
  assign n692 = ~n687 & ~n691;
  assign n685 = x46 ^ x45;
  assign n686 = x0 & n685;
  assign n693 = n692 ^ n686;
  assign n701 = n700 ^ n693;
  assign n709 = n708 ^ n701;
  assign n755 = n754 ^ n709;
  assign n759 = n758 ^ n755;
  assign n763 = n762 ^ n759;
  assign n767 = n766 ^ n763;
  assign n866 = n766 ^ n759;
  assign n867 = n763 & ~n866;
  assign n868 = n867 ^ n766;
  assign n862 = n758 ^ n754;
  assign n863 = n755 & n862;
  assign n864 = n863 ^ n709;
  assign n857 = n753 ^ n749;
  assign n858 = ~n750 & n857;
  assign n859 = n858 ^ n732;
  assign n851 = n723 ^ n716;
  assign n852 = n730 ^ n716;
  assign n853 = n851 & ~n852;
  assign n854 = n853 ^ n723;
  assign n842 = ~x11 & n159;
  assign n843 = ~x10 & n163;
  assign n844 = ~n842 & ~n843;
  assign n845 = x11 & n166;
  assign n846 = x10 & n168;
  assign n847 = ~n845 & ~n846;
  assign n848 = n844 & n847;
  assign n835 = ~x7 & n344;
  assign n836 = ~x6 & n348;
  assign n837 = ~n835 & ~n836;
  assign n838 = x7 & n351;
  assign n839 = x6 & n353;
  assign n840 = ~n838 & ~n839;
  assign n841 = n837 & n840;
  assign n849 = n848 ^ n841;
  assign n828 = x5 & n453;
  assign n829 = x4 & n457;
  assign n830 = ~n828 & ~n829;
  assign n831 = ~x5 & n460;
  assign n832 = ~x4 & n462;
  assign n833 = ~n831 & ~n832;
  assign n834 = n830 & n833;
  assign n850 = n849 ^ n834;
  assign n855 = n854 ^ n850;
  assign n813 = ~x47 & n685;
  assign n814 = x1 & n813;
  assign n815 = x47 ^ x46;
  assign n816 = ~n685 & n815;
  assign n817 = ~x47 & n816;
  assign n818 = x0 & n817;
  assign n819 = ~n814 & ~n818;
  assign n820 = x47 & n685;
  assign n821 = ~x1 & n820;
  assign n822 = x47 & n816;
  assign n823 = ~x0 & n822;
  assign n824 = ~n821 & ~n823;
  assign n825 = n819 & n824;
  assign n806 = ~x13 & n89;
  assign n807 = ~x12 & n93;
  assign n808 = ~n806 & ~n807;
  assign n809 = x13 & n96;
  assign n810 = x12 & n98;
  assign n811 = ~n809 & ~n810;
  assign n812 = n808 & n811;
  assign n826 = n825 ^ n812;
  assign n799 = x9 & n232;
  assign n800 = x8 & n234;
  assign n801 = ~n799 & ~n800;
  assign n802 = ~x9 & n225;
  assign n803 = ~x8 & n229;
  assign n804 = ~n802 & ~n803;
  assign n805 = n801 & n804;
  assign n827 = n826 ^ n805;
  assign n856 = n855 ^ n827;
  assign n860 = n859 ^ n856;
  assign n795 = n704 ^ n701;
  assign n796 = ~n708 & ~n795;
  assign n797 = n796 ^ n701;
  assign n791 = n747 ^ n733;
  assign n792 = n748 & n791;
  assign n793 = n792 ^ n740;
  assign n787 = n700 ^ n692;
  assign n788 = ~n693 & ~n787;
  assign n789 = n788 ^ n686;
  assign n779 = ~x14 & n67;
  assign n780 = n69 ^ x15;
  assign n781 = n780 ^ n69;
  assign n782 = n71 & n781;
  assign n783 = n782 ^ n69;
  assign n784 = ~n779 & ~n783;
  assign n775 = x45 ^ x0;
  assign n776 = ~n685 & n775;
  assign n777 = n776 ^ x0;
  assign n778 = x47 & ~n777;
  assign n785 = n784 ^ n778;
  assign n768 = ~x3 & n618;
  assign n769 = ~x2 & n622;
  assign n770 = ~n768 & ~n769;
  assign n771 = x3 & n625;
  assign n772 = x2 & n627;
  assign n773 = ~n771 & ~n772;
  assign n774 = n770 & n773;
  assign n786 = n785 ^ n774;
  assign n790 = n789 ^ n786;
  assign n794 = n793 ^ n790;
  assign n798 = n797 ^ n794;
  assign n861 = n860 ^ n798;
  assign n865 = n864 ^ n861;
  assign n869 = n868 ^ n865;
  assign n964 = n868 ^ n861;
  assign n965 = n865 & ~n964;
  assign n966 = n965 ^ n868;
  assign n959 = n856 ^ n798;
  assign n960 = n859 ^ n798;
  assign n961 = n959 & ~n960;
  assign n962 = n961 ^ n856;
  assign n954 = n797 ^ n793;
  assign n955 = ~n794 & n954;
  assign n956 = n955 ^ n790;
  assign n943 = ~x6 & n460;
  assign n944 = ~x5 & n462;
  assign n945 = ~n943 & ~n944;
  assign n946 = x6 & n453;
  assign n947 = x5 & n457;
  assign n948 = ~n946 & ~n947;
  assign n949 = n945 & n948;
  assign n936 = x12 & n166;
  assign n937 = x11 & n168;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~x12 & n159;
  assign n940 = ~x11 & n163;
  assign n941 = ~n939 & ~n940;
  assign n942 = n938 & n941;
  assign n950 = n949 ^ n942;
  assign n929 = x4 & n625;
  assign n930 = x3 & n627;
  assign n931 = ~n929 & ~n930;
  assign n932 = ~x4 & n618;
  assign n933 = ~x3 & n622;
  assign n934 = ~n932 & ~n933;
  assign n935 = n931 & n934;
  assign n951 = n950 ^ n935;
  assign n921 = ~x14 & n89;
  assign n922 = ~x13 & n93;
  assign n923 = ~n921 & ~n922;
  assign n924 = x14 & n96;
  assign n925 = x13 & n98;
  assign n926 = ~n924 & ~n925;
  assign n927 = n923 & n926;
  assign n914 = ~x15 & n67;
  assign n915 = n69 ^ x16;
  assign n916 = n915 ^ n69;
  assign n917 = n71 & n916;
  assign n918 = n917 ^ n69;
  assign n919 = ~n914 & ~n918;
  assign n912 = x48 ^ x47;
  assign n913 = x0 & n912;
  assign n920 = n919 ^ n913;
  assign n928 = n927 ^ n920;
  assign n952 = n951 ^ n928;
  assign n903 = x10 & n232;
  assign n904 = x9 & n234;
  assign n905 = ~n903 & ~n904;
  assign n906 = ~x10 & n225;
  assign n907 = ~x9 & n229;
  assign n908 = ~n906 & ~n907;
  assign n909 = n905 & n908;
  assign n896 = ~x2 & n820;
  assign n897 = ~x1 & n822;
  assign n898 = ~n896 & ~n897;
  assign n899 = x2 & n813;
  assign n900 = x1 & n817;
  assign n901 = ~n899 & ~n900;
  assign n902 = n898 & n901;
  assign n910 = n909 ^ n902;
  assign n889 = x8 & n351;
  assign n890 = x7 & n353;
  assign n891 = ~n889 & ~n890;
  assign n892 = ~x8 & n344;
  assign n893 = ~x7 & n348;
  assign n894 = ~n892 & ~n893;
  assign n895 = n891 & n894;
  assign n911 = n910 ^ n895;
  assign n953 = n952 ^ n911;
  assign n957 = n956 ^ n953;
  assign n884 = n850 ^ n827;
  assign n885 = n854 ^ n827;
  assign n886 = n884 & ~n885;
  assign n887 = n886 ^ n850;
  assign n880 = n789 ^ n785;
  assign n881 = n786 & n880;
  assign n882 = n881 ^ n774;
  assign n875 = n841 ^ n834;
  assign n876 = n848 ^ n834;
  assign n877 = n875 & ~n876;
  assign n878 = n877 ^ n841;
  assign n871 = n825 ^ n805;
  assign n872 = n826 & ~n871;
  assign n873 = n872 ^ n812;
  assign n870 = n778 & ~n784;
  assign n874 = n873 ^ n870;
  assign n879 = n878 ^ n874;
  assign n883 = n882 ^ n879;
  assign n888 = n887 ^ n883;
  assign n958 = n957 ^ n888;
  assign n963 = n962 ^ n958;
  assign n967 = n966 ^ n963;
  assign n1078 = n966 ^ n958;
  assign n1079 = n963 & n1078;
  assign n1080 = n1079 ^ n966;
  assign n1073 = n953 ^ n888;
  assign n1074 = n956 ^ n888;
  assign n1075 = n1073 & ~n1074;
  assign n1076 = n1075 ^ n953;
  assign n1068 = n887 ^ n882;
  assign n1069 = ~n883 & ~n1068;
  assign n1070 = n1069 ^ n879;
  assign n1057 = ~x11 & n225;
  assign n1058 = ~x10 & n229;
  assign n1059 = ~n1057 & ~n1058;
  assign n1060 = x11 & n232;
  assign n1061 = x10 & n234;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n1059 & n1062;
  assign n1050 = ~x3 & n820;
  assign n1051 = ~x2 & n822;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = x3 & n813;
  assign n1054 = x2 & n817;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1052 & n1055;
  assign n1064 = n1063 ^ n1056;
  assign n1037 = x49 & n912;
  assign n1038 = ~x1 & n1037;
  assign n1039 = x49 ^ x48;
  assign n1040 = ~n912 & n1039;
  assign n1041 = x49 & n1040;
  assign n1042 = ~x0 & n1041;
  assign n1043 = ~n1038 & ~n1042;
  assign n1044 = ~x49 & n912;
  assign n1045 = x1 & n1044;
  assign n1046 = ~x49 & n1040;
  assign n1047 = x0 & n1046;
  assign n1048 = ~n1045 & ~n1047;
  assign n1049 = n1043 & n1048;
  assign n1065 = n1064 ^ n1049;
  assign n1028 = x9 & n351;
  assign n1029 = x8 & n353;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~x9 & n344;
  assign n1032 = ~x8 & n348;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = n1030 & n1033;
  assign n1021 = x15 & n96;
  assign n1022 = x14 & n98;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~x15 & n89;
  assign n1025 = ~x14 & n93;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = n1023 & n1026;
  assign n1035 = n1034 ^ n1027;
  assign n1014 = ~x13 & n159;
  assign n1015 = ~x12 & n163;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = x13 & n166;
  assign n1018 = x12 & n168;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n1016 & n1019;
  assign n1036 = n1035 ^ n1020;
  assign n1066 = n1065 ^ n1036;
  assign n1005 = ~x7 & n460;
  assign n1006 = ~x6 & n462;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = x7 & n453;
  assign n1009 = x6 & n457;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = n1007 & n1010;
  assign n998 = x5 & n625;
  assign n999 = x4 & n627;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = ~x5 & n618;
  assign n1002 = ~x4 & n622;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = n1000 & n1003;
  assign n1012 = n1011 ^ n1004;
  assign n991 = ~x16 & n67;
  assign n992 = n69 ^ x17;
  assign n993 = n992 ^ n69;
  assign n994 = n71 & n993;
  assign n995 = n994 ^ n69;
  assign n996 = ~n991 & ~n995;
  assign n987 = x47 ^ x0;
  assign n988 = ~n912 & n987;
  assign n989 = n988 ^ x0;
  assign n990 = x49 & ~n989;
  assign n997 = n996 ^ n990;
  assign n1013 = n1012 ^ n997;
  assign n1067 = n1066 ^ n1013;
  assign n1071 = n1070 ^ n1067;
  assign n983 = n951 ^ n911;
  assign n984 = ~n952 & ~n983;
  assign n985 = n984 ^ n928;
  assign n979 = n878 ^ n873;
  assign n980 = ~n874 & ~n979;
  assign n981 = n980 ^ n870;
  assign n975 = n909 ^ n895;
  assign n976 = n910 & ~n975;
  assign n977 = n976 ^ n902;
  assign n971 = n942 ^ n935;
  assign n972 = ~n950 & n971;
  assign n973 = n972 ^ n935;
  assign n968 = n927 ^ n919;
  assign n969 = ~n920 & ~n968;
  assign n970 = n969 ^ n913;
  assign n974 = n973 ^ n970;
  assign n978 = n977 ^ n974;
  assign n982 = n981 ^ n978;
  assign n986 = n985 ^ n982;
  assign n1072 = n1071 ^ n986;
  assign n1077 = n1076 ^ n1072;
  assign n1081 = n1080 ^ n1077;
  assign n1186 = n1080 ^ n1072;
  assign n1187 = n1077 & ~n1186;
  assign n1188 = n1187 ^ n1080;
  assign n1181 = n1067 ^ n986;
  assign n1182 = n1070 ^ n986;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = n1183 ^ n1067;
  assign n1176 = n985 ^ n978;
  assign n1177 = ~n982 & n1176;
  assign n1178 = n1177 ^ n985;
  assign n1171 = n1011 ^ n997;
  assign n1172 = n1012 & ~n1171;
  assign n1173 = n1172 ^ n1004;
  assign n1162 = x2 & n1044;
  assign n1163 = x1 & n1046;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = ~x2 & n1037;
  assign n1166 = ~x1 & n1041;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = n1164 & n1167;
  assign n1155 = x4 & n813;
  assign n1156 = x3 & n817;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~x4 & n820;
  assign n1159 = ~x3 & n822;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = n1157 & n1160;
  assign n1169 = n1168 ^ n1161;
  assign n1148 = ~x16 & n89;
  assign n1149 = ~x15 & n93;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = x16 & n96;
  assign n1152 = x15 & n98;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1150 & n1153;
  assign n1170 = n1169 ^ n1154;
  assign n1174 = n1173 ^ n1170;
  assign n1144 = n1056 ^ n1049;
  assign n1145 = ~n1064 & n1144;
  assign n1146 = n1145 ^ n1049;
  assign n1142 = n990 & ~n996;
  assign n1135 = x6 & n625;
  assign n1136 = x5 & n627;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = ~x6 & n618;
  assign n1139 = ~x5 & n622;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = n1137 & n1140;
  assign n1143 = n1142 ^ n1141;
  assign n1147 = n1146 ^ n1143;
  assign n1175 = n1174 ^ n1147;
  assign n1179 = n1178 ^ n1175;
  assign n1130 = n977 ^ n973;
  assign n1131 = ~n974 & ~n1130;
  assign n1132 = n1131 ^ n970;
  assign n1127 = n1036 ^ n1013;
  assign n1128 = ~n1066 & n1127;
  assign n1129 = n1128 ^ n1013;
  assign n1133 = n1132 ^ n1129;
  assign n1122 = n1034 ^ n1020;
  assign n1123 = n1035 & ~n1122;
  assign n1124 = n1123 ^ n1027;
  assign n1113 = ~x14 & n159;
  assign n1114 = ~x13 & n163;
  assign n1115 = ~n1113 & ~n1114;
  assign n1116 = x14 & n166;
  assign n1117 = x13 & n168;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = n1115 & n1118;
  assign n1106 = ~x10 & n344;
  assign n1107 = ~x9 & n348;
  assign n1108 = ~n1106 & ~n1107;
  assign n1109 = x10 & n351;
  assign n1110 = x9 & n353;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n1108 & n1111;
  assign n1120 = n1119 ^ n1112;
  assign n1099 = ~x8 & n460;
  assign n1100 = ~x7 & n462;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = x8 & n453;
  assign n1103 = x7 & n457;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = n1101 & n1104;
  assign n1121 = n1120 ^ n1105;
  assign n1125 = n1124 ^ n1121;
  assign n1091 = ~x12 & n225;
  assign n1092 = ~x11 & n229;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = x12 & n232;
  assign n1095 = x11 & n234;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = n1093 & n1096;
  assign n1084 = ~x17 & n67;
  assign n1085 = n69 ^ x18;
  assign n1086 = n1085 ^ n69;
  assign n1087 = n71 & n1086;
  assign n1088 = n1087 ^ n69;
  assign n1089 = ~n1084 & ~n1088;
  assign n1082 = x50 ^ x49;
  assign n1083 = x0 & n1082;
  assign n1090 = n1089 ^ n1083;
  assign n1098 = n1097 ^ n1090;
  assign n1126 = n1125 ^ n1098;
  assign n1134 = n1133 ^ n1126;
  assign n1180 = n1179 ^ n1134;
  assign n1185 = n1184 ^ n1180;
  assign n1189 = n1188 ^ n1185;
  assign n1312 = n1188 ^ n1180;
  assign n1313 = ~n1185 & ~n1312;
  assign n1314 = n1313 ^ n1188;
  assign n1307 = n1175 ^ n1134;
  assign n1308 = n1178 ^ n1134;
  assign n1309 = ~n1307 & n1308;
  assign n1310 = n1309 ^ n1175;
  assign n1302 = n1129 ^ n1126;
  assign n1303 = n1133 & ~n1302;
  assign n1304 = n1303 ^ n1126;
  assign n1297 = n1146 ^ n1142;
  assign n1298 = ~n1143 & n1297;
  assign n1299 = n1298 ^ n1141;
  assign n1288 = x17 & n96;
  assign n1289 = x16 & n98;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~x17 & n89;
  assign n1292 = ~x16 & n93;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n1290 & n1293;
  assign n1275 = ~x51 & n1082;
  assign n1276 = x1 & n1275;
  assign n1277 = x51 ^ x50;
  assign n1278 = ~n1082 & n1277;
  assign n1279 = ~x51 & n1278;
  assign n1280 = x0 & n1279;
  assign n1281 = ~n1276 & ~n1280;
  assign n1282 = x51 & n1082;
  assign n1283 = ~x1 & n1282;
  assign n1284 = x51 & n1278;
  assign n1285 = ~x0 & n1284;
  assign n1286 = ~n1283 & ~n1285;
  assign n1287 = n1281 & n1286;
  assign n1295 = n1294 ^ n1287;
  assign n1268 = x11 & n351;
  assign n1269 = x10 & n353;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~x11 & n344;
  assign n1272 = ~x10 & n348;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = n1270 & n1273;
  assign n1296 = n1295 ^ n1274;
  assign n1300 = n1299 ^ n1296;
  assign n1264 = n1161 ^ n1154;
  assign n1265 = ~n1169 & n1264;
  assign n1266 = n1265 ^ n1154;
  assign n1260 = n1097 ^ n1089;
  assign n1261 = ~n1090 & ~n1260;
  assign n1262 = n1261 ^ n1083;
  assign n1253 = ~x18 & n67;
  assign n1254 = n69 ^ x19;
  assign n1255 = n1254 ^ n69;
  assign n1256 = n71 & n1255;
  assign n1257 = n1256 ^ n69;
  assign n1258 = ~n1253 & ~n1257;
  assign n1249 = x49 ^ x0;
  assign n1250 = ~n1082 & n1249;
  assign n1251 = n1250 ^ x0;
  assign n1252 = x51 & ~n1251;
  assign n1259 = n1258 ^ n1252;
  assign n1263 = n1262 ^ n1259;
  assign n1267 = n1266 ^ n1263;
  assign n1301 = n1300 ^ n1267;
  assign n1305 = n1304 ^ n1301;
  assign n1245 = n1173 ^ n1147;
  assign n1246 = n1174 & n1245;
  assign n1247 = n1246 ^ n1170;
  assign n1241 = n1121 ^ n1098;
  assign n1242 = ~n1125 & ~n1241;
  assign n1243 = n1242 ^ n1098;
  assign n1236 = n1112 ^ n1105;
  assign n1237 = ~n1120 & n1236;
  assign n1238 = n1237 ^ n1105;
  assign n1227 = ~x9 & n460;
  assign n1228 = ~x8 & n462;
  assign n1229 = ~n1227 & ~n1228;
  assign n1230 = x9 & n453;
  assign n1231 = x8 & n457;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = n1229 & n1232;
  assign n1220 = ~x15 & n159;
  assign n1221 = ~x14 & n163;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = x15 & n166;
  assign n1224 = x14 & n168;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = n1222 & n1225;
  assign n1234 = n1233 ^ n1226;
  assign n1213 = ~x7 & n618;
  assign n1214 = ~x6 & n622;
  assign n1215 = ~n1213 & ~n1214;
  assign n1216 = x7 & n625;
  assign n1217 = x6 & n627;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n1215 & n1218;
  assign n1235 = n1234 ^ n1219;
  assign n1239 = n1238 ^ n1235;
  assign n1204 = x5 & n813;
  assign n1205 = x4 & n817;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = ~x5 & n820;
  assign n1208 = ~x4 & n822;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n1206 & n1209;
  assign n1197 = x13 & n232;
  assign n1198 = x12 & n234;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~x13 & n225;
  assign n1201 = ~x12 & n229;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = n1199 & n1202;
  assign n1211 = n1210 ^ n1203;
  assign n1190 = ~x3 & n1037;
  assign n1191 = ~x2 & n1041;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = x3 & n1044;
  assign n1194 = x2 & n1046;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1192 & n1195;
  assign n1212 = n1211 ^ n1196;
  assign n1240 = n1239 ^ n1212;
  assign n1244 = n1243 ^ n1240;
  assign n1248 = n1247 ^ n1244;
  assign n1306 = n1305 ^ n1248;
  assign n1311 = n1310 ^ n1306;
  assign n1315 = n1314 ^ n1311;
  assign n1435 = n1314 ^ n1306;
  assign n1436 = ~n1311 & n1435;
  assign n1437 = n1436 ^ n1314;
  assign n1430 = n1301 ^ n1248;
  assign n1431 = n1304 ^ n1248;
  assign n1432 = n1430 & ~n1431;
  assign n1433 = n1432 ^ n1301;
  assign n1424 = n1247 ^ n1240;
  assign n1425 = n1247 ^ n1243;
  assign n1426 = n1424 & n1425;
  assign n1427 = n1426 ^ n1240;
  assign n1420 = n1296 ^ n1267;
  assign n1421 = n1299 ^ n1267;
  assign n1422 = ~n1420 & n1421;
  assign n1423 = n1422 ^ n1296;
  assign n1428 = n1427 ^ n1423;
  assign n1414 = n1235 ^ n1212;
  assign n1415 = n1238 ^ n1212;
  assign n1416 = n1414 & ~n1415;
  assign n1417 = n1416 ^ n1235;
  assign n1410 = n1266 ^ n1262;
  assign n1411 = ~n1263 & n1410;
  assign n1412 = n1411 ^ n1259;
  assign n1401 = ~x8 & n618;
  assign n1402 = ~x7 & n622;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = x8 & n625;
  assign n1405 = x7 & n627;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = n1403 & n1406;
  assign n1394 = ~x10 & n460;
  assign n1395 = ~x9 & n462;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = x10 & n453;
  assign n1398 = x9 & n457;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = n1396 & n1399;
  assign n1408 = n1407 ^ n1400;
  assign n1393 = n1252 & ~n1258;
  assign n1409 = n1408 ^ n1393;
  assign n1413 = n1412 ^ n1409;
  assign n1418 = n1417 ^ n1413;
  assign n1388 = n1287 ^ n1274;
  assign n1389 = ~n1295 & n1388;
  assign n1390 = n1389 ^ n1274;
  assign n1384 = n1210 ^ n1196;
  assign n1385 = n1211 & ~n1384;
  assign n1386 = n1385 ^ n1203;
  assign n1381 = n1233 ^ n1219;
  assign n1382 = n1234 & ~n1381;
  assign n1383 = n1382 ^ n1226;
  assign n1387 = n1386 ^ n1383;
  assign n1391 = n1390 ^ n1387;
  assign n1370 = ~x6 & n820;
  assign n1371 = ~x5 & n822;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = x6 & n813;
  assign n1374 = x5 & n817;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = n1372 & n1375;
  assign n1363 = ~x4 & n1037;
  assign n1364 = ~x3 & n1041;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = x4 & n1044;
  assign n1367 = x3 & n1046;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n1365 & n1368;
  assign n1377 = n1376 ^ n1369;
  assign n1356 = ~x18 & n89;
  assign n1357 = ~x17 & n93;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = x18 & n96;
  assign n1360 = x17 & n98;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = n1358 & n1361;
  assign n1378 = n1377 ^ n1362;
  assign n1348 = ~x14 & n225;
  assign n1349 = ~x13 & n229;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = x14 & n232;
  assign n1352 = x13 & n234;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = n1350 & n1353;
  assign n1341 = ~x19 & n67;
  assign n1342 = n69 ^ x20;
  assign n1343 = n1342 ^ n69;
  assign n1344 = n71 & n1343;
  assign n1345 = n1344 ^ n69;
  assign n1346 = ~n1341 & ~n1345;
  assign n1339 = x52 ^ x51;
  assign n1340 = x0 & n1339;
  assign n1347 = n1346 ^ n1340;
  assign n1355 = n1354 ^ n1347;
  assign n1379 = n1378 ^ n1355;
  assign n1330 = ~x12 & n344;
  assign n1331 = ~x11 & n348;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = x12 & n351;
  assign n1334 = x11 & n353;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = n1332 & n1335;
  assign n1323 = ~x2 & n1282;
  assign n1324 = ~x1 & n1284;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = x2 & n1275;
  assign n1327 = x1 & n1279;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = n1325 & n1328;
  assign n1337 = n1336 ^ n1329;
  assign n1316 = x16 & n166;
  assign n1317 = x15 & n168;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~x16 & n159;
  assign n1320 = ~x15 & n163;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = n1318 & n1321;
  assign n1338 = n1337 ^ n1322;
  assign n1380 = n1379 ^ n1338;
  assign n1392 = n1391 ^ n1380;
  assign n1419 = n1418 ^ n1392;
  assign n1429 = n1428 ^ n1419;
  assign n1434 = n1433 ^ n1429;
  assign n1438 = n1437 ^ n1434;
  assign n1574 = n1437 ^ n1429;
  assign n1575 = n1434 & ~n1574;
  assign n1576 = n1575 ^ n1437;
  assign n1570 = n1423 ^ n1419;
  assign n1571 = ~n1428 & n1570;
  assign n1572 = n1571 ^ n1419;
  assign n1566 = n1418 ^ n1391;
  assign n1567 = ~n1392 & n1566;
  assign n1568 = n1567 ^ n1380;
  assign n1561 = n1417 ^ n1409;
  assign n1562 = n1417 ^ n1412;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = n1563 ^ n1409;
  assign n1555 = n1390 ^ n1386;
  assign n1556 = n1387 & ~n1555;
  assign n1557 = n1556 ^ n1383;
  assign n1550 = n1369 ^ n1362;
  assign n1551 = n1376 ^ n1362;
  assign n1552 = n1550 & ~n1551;
  assign n1553 = n1552 ^ n1369;
  assign n1541 = x19 & n96;
  assign n1542 = x18 & n98;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = ~x19 & n89;
  assign n1545 = ~x18 & n93;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = n1543 & n1546;
  assign n1537 = x51 ^ x0;
  assign n1538 = ~n1339 & n1537;
  assign n1539 = n1538 ^ x0;
  assign n1540 = x53 & ~n1539;
  assign n1548 = n1547 ^ n1540;
  assign n1530 = x9 & n625;
  assign n1531 = x8 & n627;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = ~x9 & n618;
  assign n1534 = ~x8 & n622;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = n1532 & n1535;
  assign n1549 = n1548 ^ n1536;
  assign n1554 = n1553 ^ n1549;
  assign n1558 = n1557 ^ n1554;
  assign n1525 = n1336 ^ n1322;
  assign n1526 = n1337 & ~n1525;
  assign n1527 = n1526 ^ n1329;
  assign n1522 = n1354 ^ n1346;
  assign n1523 = ~n1347 & ~n1522;
  assign n1524 = n1523 ^ n1340;
  assign n1528 = n1527 ^ n1524;
  assign n1514 = ~x20 & n67;
  assign n1515 = n69 ^ x21;
  assign n1516 = n1515 ^ n69;
  assign n1517 = n71 & n1516;
  assign n1518 = n1517 ^ n69;
  assign n1519 = ~n1514 & ~n1518;
  assign n1507 = ~x17 & n159;
  assign n1508 = ~x16 & n163;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = x17 & n166;
  assign n1511 = x16 & n168;
  assign n1512 = ~n1510 & ~n1511;
  assign n1513 = n1509 & n1512;
  assign n1520 = n1519 ^ n1513;
  assign n1500 = ~x11 & n460;
  assign n1501 = ~x10 & n462;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = x11 & n453;
  assign n1504 = x10 & n457;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = n1502 & n1505;
  assign n1521 = n1520 ^ n1506;
  assign n1529 = n1528 ^ n1521;
  assign n1559 = n1558 ^ n1529;
  assign n1496 = n1378 ^ n1338;
  assign n1497 = ~n1379 & ~n1496;
  assign n1498 = n1497 ^ n1355;
  assign n1492 = n1407 ^ n1393;
  assign n1493 = n1408 & n1492;
  assign n1494 = n1493 ^ n1400;
  assign n1482 = ~x15 & n225;
  assign n1483 = ~x14 & n229;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = x15 & n232;
  assign n1486 = x14 & n234;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = n1484 & n1487;
  assign n1475 = x7 & n813;
  assign n1476 = x6 & n817;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = ~x7 & n820;
  assign n1479 = ~x6 & n822;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = n1477 & n1480;
  assign n1489 = n1488 ^ n1481;
  assign n1468 = ~x5 & n1037;
  assign n1469 = ~x4 & n1041;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = x5 & n1044;
  assign n1472 = x4 & n1046;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = n1470 & n1473;
  assign n1490 = n1489 ^ n1474;
  assign n1459 = x3 & n1275;
  assign n1460 = x2 & n1279;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~x3 & n1282;
  assign n1463 = ~x2 & n1284;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = n1461 & n1464;
  assign n1452 = ~x13 & n344;
  assign n1453 = ~x12 & n348;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = x13 & n351;
  assign n1456 = x12 & n353;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = n1454 & n1457;
  assign n1466 = n1465 ^ n1458;
  assign n1439 = x53 & n1339;
  assign n1440 = ~x1 & n1439;
  assign n1441 = x53 ^ x52;
  assign n1442 = ~n1339 & n1441;
  assign n1443 = x53 & n1442;
  assign n1444 = ~x0 & n1443;
  assign n1445 = ~n1440 & ~n1444;
  assign n1446 = ~x53 & n1339;
  assign n1447 = x1 & n1446;
  assign n1448 = ~x53 & n1442;
  assign n1449 = x0 & n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = n1445 & n1450;
  assign n1467 = n1466 ^ n1451;
  assign n1491 = n1490 ^ n1467;
  assign n1495 = n1494 ^ n1491;
  assign n1499 = n1498 ^ n1495;
  assign n1560 = n1559 ^ n1499;
  assign n1565 = n1564 ^ n1560;
  assign n1569 = n1568 ^ n1565;
  assign n1573 = n1572 ^ n1569;
  assign n1577 = n1576 ^ n1573;
  assign n1707 = n1576 ^ n1569;
  assign n1708 = ~n1573 & ~n1707;
  assign n1709 = n1708 ^ n1576;
  assign n1702 = n1568 ^ n1560;
  assign n1703 = n1568 ^ n1564;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = n1704 ^ n1560;
  assign n1698 = n1559 ^ n1495;
  assign n1699 = ~n1499 & n1698;
  assign n1700 = n1699 ^ n1498;
  assign n1692 = n1554 ^ n1529;
  assign n1693 = n1557 ^ n1529;
  assign n1694 = ~n1692 & n1693;
  assign n1695 = n1694 ^ n1554;
  assign n1687 = n1553 ^ n1548;
  assign n1688 = n1549 & ~n1687;
  assign n1689 = n1688 ^ n1536;
  assign n1679 = ~x21 & n67;
  assign n1680 = n69 ^ x22;
  assign n1681 = n1680 ^ n69;
  assign n1682 = n71 & n1681;
  assign n1683 = n1682 ^ n69;
  assign n1684 = ~n1679 & ~n1683;
  assign n1671 = x2 & n1446;
  assign n1672 = x1 & n1448;
  assign n1673 = ~n1671 & ~n1672;
  assign n1674 = ~x2 & n1439;
  assign n1675 = ~x1 & n1443;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = n1673 & n1676;
  assign n1664 = x4 & n1275;
  assign n1665 = x3 & n1279;
  assign n1666 = ~n1664 & ~n1665;
  assign n1667 = ~x4 & n1282;
  assign n1668 = ~x3 & n1284;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n1666 & n1669;
  assign n1678 = n1677 ^ n1670;
  assign n1685 = n1684 ^ n1678;
  assign n1655 = x20 & n96;
  assign n1656 = x19 & n98;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = ~x20 & n89;
  assign n1659 = ~x19 & n93;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = n1657 & n1660;
  assign n1653 = x54 ^ x53;
  assign n1654 = x0 & n1653;
  assign n1662 = n1661 ^ n1654;
  assign n1646 = ~x16 & n225;
  assign n1647 = ~x15 & n229;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = x16 & n232;
  assign n1650 = x15 & n234;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = n1648 & n1651;
  assign n1663 = n1662 ^ n1652;
  assign n1686 = n1685 ^ n1663;
  assign n1690 = n1689 ^ n1686;
  assign n1641 = n1488 ^ n1474;
  assign n1642 = n1489 & ~n1641;
  assign n1643 = n1642 ^ n1481;
  assign n1632 = ~x12 & n460;
  assign n1633 = ~x11 & n462;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = x12 & n453;
  assign n1636 = x11 & n457;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n1634 & n1637;
  assign n1625 = ~x18 & n159;
  assign n1626 = ~x17 & n163;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = x18 & n166;
  assign n1629 = x17 & n168;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1627 & n1630;
  assign n1639 = n1638 ^ n1631;
  assign n1618 = ~x10 & n618;
  assign n1619 = ~x9 & n622;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = x10 & n625;
  assign n1622 = x9 & n627;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = n1620 & n1623;
  assign n1640 = n1639 ^ n1624;
  assign n1644 = n1643 ^ n1640;
  assign n1609 = ~x6 & n1037;
  assign n1610 = ~x5 & n1041;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = x6 & n1044;
  assign n1613 = x5 & n1046;
  assign n1614 = ~n1612 & ~n1613;
  assign n1615 = n1611 & n1614;
  assign n1602 = x8 & n813;
  assign n1603 = x7 & n817;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = ~x8 & n820;
  assign n1606 = ~x7 & n822;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n1604 & n1607;
  assign n1616 = n1615 ^ n1608;
  assign n1595 = x14 & n351;
  assign n1596 = x13 & n353;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~x14 & n344;
  assign n1599 = ~x13 & n348;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = n1597 & n1600;
  assign n1617 = n1616 ^ n1601;
  assign n1645 = n1644 ^ n1617;
  assign n1691 = n1690 ^ n1645;
  assign n1696 = n1695 ^ n1691;
  assign n1591 = n1494 ^ n1490;
  assign n1592 = n1491 & ~n1591;
  assign n1593 = n1592 ^ n1467;
  assign n1587 = n1524 ^ n1521;
  assign n1588 = n1528 & ~n1587;
  assign n1589 = n1588 ^ n1521;
  assign n1583 = n1458 ^ n1451;
  assign n1584 = ~n1466 & n1583;
  assign n1585 = n1584 ^ n1451;
  assign n1579 = n1513 ^ n1506;
  assign n1580 = n1520 & ~n1579;
  assign n1581 = n1580 ^ n1519;
  assign n1578 = n1540 & ~n1547;
  assign n1582 = n1581 ^ n1578;
  assign n1586 = n1585 ^ n1582;
  assign n1590 = n1589 ^ n1586;
  assign n1594 = n1593 ^ n1590;
  assign n1697 = n1696 ^ n1594;
  assign n1701 = n1700 ^ n1697;
  assign n1706 = n1705 ^ n1701;
  assign n1710 = n1709 ^ n1706;
  assign n1858 = n1709 ^ n1701;
  assign n1859 = n1706 & n1858;
  assign n1860 = n1859 ^ n1709;
  assign n1854 = n1700 ^ n1696;
  assign n1855 = n1697 & ~n1854;
  assign n1856 = n1855 ^ n1594;
  assign n1849 = n1695 ^ n1690;
  assign n1850 = ~n1691 & n1849;
  assign n1851 = n1850 ^ n1645;
  assign n1846 = n1593 ^ n1589;
  assign n1847 = ~n1590 & ~n1846;
  assign n1848 = n1847 ^ n1586;
  assign n1852 = n1851 ^ n1848;
  assign n1841 = n1689 ^ n1685;
  assign n1842 = ~n1686 & ~n1841;
  assign n1843 = n1842 ^ n1663;
  assign n1837 = n1585 ^ n1581;
  assign n1838 = ~n1582 & ~n1837;
  assign n1839 = n1838 ^ n1578;
  assign n1827 = x9 & n813;
  assign n1828 = x8 & n817;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~x9 & n820;
  assign n1831 = ~x8 & n822;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1829 & n1832;
  assign n1820 = ~x17 & n225;
  assign n1821 = ~x16 & n229;
  assign n1822 = ~n1820 & ~n1821;
  assign n1823 = x17 & n232;
  assign n1824 = x16 & n234;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = n1822 & n1825;
  assign n1834 = n1833 ^ n1826;
  assign n1813 = ~x7 & n1037;
  assign n1814 = ~x6 & n1041;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = x7 & n1044;
  assign n1817 = x6 & n1046;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = n1815 & n1818;
  assign n1835 = n1834 ^ n1819;
  assign n1804 = ~x21 & n89;
  assign n1805 = ~x20 & n93;
  assign n1806 = ~n1804 & ~n1805;
  assign n1807 = x21 & n96;
  assign n1808 = x20 & n98;
  assign n1809 = ~n1807 & ~n1808;
  assign n1810 = n1806 & n1809;
  assign n1800 = x53 ^ x0;
  assign n1801 = ~n1653 & n1800;
  assign n1802 = n1801 ^ x0;
  assign n1803 = x55 & ~n1802;
  assign n1811 = n1810 ^ n1803;
  assign n1792 = ~x11 & n618;
  assign n1793 = ~x10 & n622;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = x11 & n625;
  assign n1796 = x10 & n627;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = n1794 & n1797;
  assign n1785 = ~x13 & n460;
  assign n1786 = ~x12 & n462;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = x13 & n453;
  assign n1789 = x12 & n457;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = n1787 & n1790;
  assign n1799 = n1798 ^ n1791;
  assign n1812 = n1811 ^ n1799;
  assign n1836 = n1835 ^ n1812;
  assign n1840 = n1839 ^ n1836;
  assign n1844 = n1843 ^ n1840;
  assign n1779 = n1640 ^ n1617;
  assign n1780 = n1643 ^ n1617;
  assign n1781 = n1779 & ~n1780;
  assign n1782 = n1781 ^ n1640;
  assign n1774 = n1654 ^ n1652;
  assign n1775 = n1661 ^ n1652;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n1776 ^ n1654;
  assign n1770 = n1684 ^ n1670;
  assign n1771 = ~n1678 & n1770;
  assign n1772 = n1771 ^ n1684;
  assign n1767 = n1638 ^ n1624;
  assign n1768 = n1639 & ~n1767;
  assign n1769 = n1768 ^ n1631;
  assign n1773 = n1772 ^ n1769;
  assign n1778 = n1777 ^ n1773;
  assign n1783 = n1782 ^ n1778;
  assign n1762 = n1608 ^ n1601;
  assign n1763 = ~n1616 & n1762;
  assign n1764 = n1763 ^ n1601;
  assign n1754 = ~x22 & n67;
  assign n1755 = n69 ^ x23;
  assign n1756 = n1755 ^ n69;
  assign n1757 = n71 & n1756;
  assign n1758 = n1757 ^ n69;
  assign n1759 = ~n1754 & ~n1758;
  assign n1747 = x19 & n166;
  assign n1748 = x18 & n168;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~x19 & n159;
  assign n1751 = ~x18 & n163;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = n1749 & n1752;
  assign n1760 = n1759 ^ n1753;
  assign n1734 = x55 & n1653;
  assign n1735 = ~x1 & n1734;
  assign n1736 = x55 ^ x54;
  assign n1737 = ~n1653 & n1736;
  assign n1738 = x55 & n1737;
  assign n1739 = ~x0 & n1738;
  assign n1740 = ~n1735 & ~n1739;
  assign n1741 = ~x55 & n1653;
  assign n1742 = x1 & n1741;
  assign n1743 = ~x55 & n1737;
  assign n1744 = x0 & n1743;
  assign n1745 = ~n1742 & ~n1744;
  assign n1746 = n1740 & n1745;
  assign n1761 = n1760 ^ n1746;
  assign n1765 = n1764 ^ n1761;
  assign n1725 = x5 & n1275;
  assign n1726 = x4 & n1279;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = ~x5 & n1282;
  assign n1729 = ~x4 & n1284;
  assign n1730 = ~n1728 & ~n1729;
  assign n1731 = n1727 & n1730;
  assign n1718 = x15 & n351;
  assign n1719 = x14 & n353;
  assign n1720 = ~n1718 & ~n1719;
  assign n1721 = ~x15 & n344;
  assign n1722 = ~x14 & n348;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = n1720 & n1723;
  assign n1732 = n1731 ^ n1724;
  assign n1711 = ~x3 & n1439;
  assign n1712 = ~x2 & n1443;
  assign n1713 = ~n1711 & ~n1712;
  assign n1714 = x3 & n1446;
  assign n1715 = x2 & n1448;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = n1713 & n1716;
  assign n1733 = n1732 ^ n1717;
  assign n1766 = n1765 ^ n1733;
  assign n1784 = n1783 ^ n1766;
  assign n1845 = n1844 ^ n1784;
  assign n1853 = n1852 ^ n1845;
  assign n1857 = n1856 ^ n1853;
  assign n1861 = n1860 ^ n1857;
  assign n2002 = n1860 ^ n1853;
  assign n2003 = n1857 & ~n2002;
  assign n2004 = n2003 ^ n1860;
  assign n1998 = n1848 ^ n1845;
  assign n1999 = n1852 & n1998;
  assign n2000 = n1999 ^ n1845;
  assign n1993 = n1840 ^ n1784;
  assign n1994 = n1843 ^ n1784;
  assign n1995 = n1993 & ~n1994;
  assign n1996 = n1995 ^ n1840;
  assign n1988 = n1778 ^ n1766;
  assign n1989 = n1783 & ~n1988;
  assign n1990 = n1989 ^ n1766;
  assign n1984 = n1839 ^ n1835;
  assign n1985 = n1836 & n1984;
  assign n1986 = n1985 ^ n1812;
  assign n1979 = n1777 ^ n1769;
  assign n1980 = ~n1773 & ~n1979;
  assign n1981 = n1980 ^ n1777;
  assign n1976 = n1811 ^ n1798;
  assign n1977 = n1799 & ~n1976;
  assign n1978 = n1977 ^ n1791;
  assign n1982 = n1981 ^ n1978;
  assign n1972 = n1724 ^ n1717;
  assign n1973 = ~n1732 & n1972;
  assign n1974 = n1973 ^ n1717;
  assign n1970 = n1803 & ~n1810;
  assign n1963 = ~x12 & n618;
  assign n1964 = ~x11 & n622;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = x12 & n625;
  assign n1967 = x11 & n627;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = n1965 & n1968;
  assign n1971 = n1970 ^ n1969;
  assign n1975 = n1974 ^ n1971;
  assign n1983 = n1982 ^ n1975;
  assign n1987 = n1986 ^ n1983;
  assign n1991 = n1990 ^ n1987;
  assign n1958 = n1761 ^ n1733;
  assign n1959 = ~n1765 & n1958;
  assign n1960 = n1959 ^ n1733;
  assign n1953 = n1826 ^ n1819;
  assign n1954 = ~n1834 & n1953;
  assign n1955 = n1954 ^ n1819;
  assign n1950 = n1753 ^ n1746;
  assign n1951 = n1760 & ~n1950;
  assign n1952 = n1951 ^ n1759;
  assign n1956 = n1955 ^ n1952;
  assign n1941 = ~x20 & n159;
  assign n1942 = ~x19 & n163;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = x20 & n166;
  assign n1945 = x19 & n168;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = n1943 & n1946;
  assign n1934 = ~x2 & n1734;
  assign n1935 = ~x1 & n1738;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = x2 & n1741;
  assign n1938 = x1 & n1743;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = n1936 & n1939;
  assign n1948 = n1947 ^ n1940;
  assign n1927 = ~x14 & n460;
  assign n1928 = ~x13 & n462;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = x14 & n453;
  assign n1931 = x13 & n457;
  assign n1932 = ~n1930 & ~n1931;
  assign n1933 = n1929 & n1932;
  assign n1949 = n1948 ^ n1933;
  assign n1957 = n1956 ^ n1949;
  assign n1961 = n1960 ^ n1957;
  assign n1918 = ~x23 & n67;
  assign n1919 = n69 ^ x24;
  assign n1920 = n1919 ^ n69;
  assign n1921 = n71 & n1920;
  assign n1922 = n1921 ^ n69;
  assign n1923 = ~n1918 & ~n1922;
  assign n1910 = ~x4 & n1439;
  assign n1911 = ~x3 & n1443;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = x4 & n1446;
  assign n1914 = x3 & n1448;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = n1912 & n1915;
  assign n1903 = ~x6 & n1282;
  assign n1904 = ~x5 & n1284;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = x6 & n1275;
  assign n1907 = x5 & n1279;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = n1905 & n1908;
  assign n1917 = n1916 ^ n1909;
  assign n1924 = n1923 ^ n1917;
  assign n1894 = ~x22 & n89;
  assign n1895 = ~x21 & n93;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = x22 & n96;
  assign n1898 = x21 & n98;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = n1896 & n1899;
  assign n1892 = x56 ^ x55;
  assign n1893 = x0 & n1892;
  assign n1901 = n1900 ^ n1893;
  assign n1885 = ~x18 & n225;
  assign n1886 = ~x17 & n229;
  assign n1887 = ~n1885 & ~n1886;
  assign n1888 = x18 & n232;
  assign n1889 = x17 & n234;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = n1887 & n1890;
  assign n1902 = n1901 ^ n1891;
  assign n1925 = n1924 ^ n1902;
  assign n1876 = x10 & n813;
  assign n1877 = x9 & n817;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~x10 & n820;
  assign n1880 = ~x9 & n822;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n1878 & n1881;
  assign n1869 = x8 & n1044;
  assign n1870 = x7 & n1046;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = ~x8 & n1037;
  assign n1873 = ~x7 & n1041;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = n1871 & n1874;
  assign n1883 = n1882 ^ n1875;
  assign n1862 = ~x16 & n344;
  assign n1863 = ~x15 & n348;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = x16 & n351;
  assign n1866 = x15 & n353;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = n1864 & n1867;
  assign n1884 = n1883 ^ n1868;
  assign n1926 = n1925 ^ n1884;
  assign n1962 = n1961 ^ n1926;
  assign n1992 = n1991 ^ n1962;
  assign n1997 = n1996 ^ n1992;
  assign n2001 = n2000 ^ n1997;
  assign n2005 = n2004 ^ n2001;
  assign n2167 = n2004 ^ n1997;
  assign n2168 = n2001 & ~n2167;
  assign n2169 = n2168 ^ n2004;
  assign n2163 = n1996 ^ n1991;
  assign n2164 = ~n1992 & n2163;
  assign n2165 = n2164 ^ n1962;
  assign n2158 = n1990 ^ n1986;
  assign n2159 = n1987 & ~n2158;
  assign n2160 = n2159 ^ n1983;
  assign n2153 = n1952 ^ n1949;
  assign n2154 = ~n1956 & n2153;
  assign n2155 = n2154 ^ n1949;
  assign n2149 = n1923 ^ n1909;
  assign n2150 = ~n1917 & n2149;
  assign n2151 = n2150 ^ n1923;
  assign n2144 = n1875 ^ n1868;
  assign n2145 = n1882 ^ n1868;
  assign n2146 = n2144 & ~n2145;
  assign n2147 = n2146 ^ n1875;
  assign n2136 = x23 & n96;
  assign n2137 = x22 & n98;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = ~x23 & n89;
  assign n2140 = ~x22 & n93;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = n2138 & n2141;
  assign n2132 = x55 ^ x0;
  assign n2133 = ~n1892 & n2132;
  assign n2134 = n2133 ^ x0;
  assign n2135 = x57 & ~n2134;
  assign n2143 = n2142 ^ n2135;
  assign n2148 = n2147 ^ n2143;
  assign n2152 = n2151 ^ n2148;
  assign n2156 = n2155 ^ n2152;
  assign n2121 = x7 & n1275;
  assign n2122 = x6 & n1279;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = ~x7 & n1282;
  assign n2125 = ~x6 & n1284;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = n2123 & n2126;
  assign n2114 = ~x17 & n344;
  assign n2115 = ~x16 & n348;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = x17 & n351;
  assign n2118 = x16 & n353;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = n2116 & n2119;
  assign n2128 = n2127 ^ n2120;
  assign n2107 = x5 & n1446;
  assign n2108 = x4 & n1448;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~x5 & n1439;
  assign n2111 = ~x4 & n1443;
  assign n2112 = ~n2110 & ~n2111;
  assign n2113 = n2109 & n2112;
  assign n2129 = n2128 ^ n2113;
  assign n2098 = ~x11 & n820;
  assign n2099 = ~x10 & n822;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = x11 & n813;
  assign n2102 = x10 & n817;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = n2100 & n2103;
  assign n2091 = ~x19 & n225;
  assign n2092 = ~x18 & n229;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = x19 & n232;
  assign n2095 = x18 & n234;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = n2093 & n2096;
  assign n2105 = n2104 ^ n2097;
  assign n2084 = ~x9 & n1037;
  assign n2085 = ~x8 & n1041;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = x9 & n1044;
  assign n2088 = x8 & n1046;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n2086 & n2089;
  assign n2106 = n2105 ^ n2090;
  assign n2130 = n2129 ^ n2106;
  assign n2076 = ~x24 & n67;
  assign n2077 = n69 ^ x25;
  assign n2078 = n2077 ^ n69;
  assign n2079 = n71 & n2078;
  assign n2080 = n2079 ^ n69;
  assign n2081 = ~n2076 & ~n2080;
  assign n2069 = x15 & n453;
  assign n2070 = x14 & n457;
  assign n2071 = ~n2069 & ~n2070;
  assign n2072 = ~x15 & n460;
  assign n2073 = ~x14 & n462;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = n2071 & n2074;
  assign n2082 = n2081 ^ n2075;
  assign n2062 = x3 & n1741;
  assign n2063 = x2 & n1743;
  assign n2064 = ~n2062 & ~n2063;
  assign n2065 = ~x3 & n1734;
  assign n2066 = ~x2 & n1738;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = n2064 & n2067;
  assign n2083 = n2082 ^ n2068;
  assign n2131 = n2130 ^ n2083;
  assign n2157 = n2156 ^ n2131;
  assign n2161 = n2160 ^ n2157;
  assign n2056 = n1978 ^ n1975;
  assign n2057 = n1981 ^ n1975;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = n2058 ^ n1978;
  assign n2053 = n1957 ^ n1926;
  assign n2054 = ~n1961 & ~n2053;
  assign n2055 = n2054 ^ n1926;
  assign n2060 = n2059 ^ n2055;
  assign n2048 = n1902 ^ n1884;
  assign n2049 = n1924 ^ n1884;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = n2050 ^ n1902;
  assign n2044 = n1974 ^ n1970;
  assign n2045 = ~n1971 & n2044;
  assign n2046 = n2045 ^ n1969;
  assign n2038 = n1940 ^ n1933;
  assign n2039 = n1947 ^ n1933;
  assign n2040 = n2038 & ~n2039;
  assign n2041 = n2040 ^ n1940;
  assign n2035 = n1900 ^ n1891;
  assign n2036 = ~n1901 & ~n2035;
  assign n2037 = n2036 ^ n1893;
  assign n2042 = n2041 ^ n2037;
  assign n2026 = ~x21 & n159;
  assign n2027 = ~x20 & n163;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = x21 & n166;
  assign n2030 = x20 & n168;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = n2028 & n2031;
  assign n2013 = x57 & n1892;
  assign n2014 = ~x1 & n2013;
  assign n2015 = x57 ^ x56;
  assign n2016 = ~n1892 & n2015;
  assign n2017 = x57 & n2016;
  assign n2018 = ~x0 & n2017;
  assign n2019 = ~n2014 & ~n2018;
  assign n2020 = ~x57 & n1892;
  assign n2021 = x1 & n2020;
  assign n2022 = ~x57 & n2016;
  assign n2023 = x0 & n2022;
  assign n2024 = ~n2021 & ~n2023;
  assign n2025 = n2019 & n2024;
  assign n2033 = n2032 ^ n2025;
  assign n2006 = ~x13 & n618;
  assign n2007 = ~x12 & n622;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = x13 & n625;
  assign n2010 = x12 & n627;
  assign n2011 = ~n2009 & ~n2010;
  assign n2012 = n2008 & n2011;
  assign n2034 = n2033 ^ n2012;
  assign n2043 = n2042 ^ n2034;
  assign n2047 = n2046 ^ n2043;
  assign n2052 = n2051 ^ n2047;
  assign n2061 = n2060 ^ n2052;
  assign n2162 = n2161 ^ n2061;
  assign n2166 = n2165 ^ n2162;
  assign n2170 = n2169 ^ n2166;
  assign n2326 = n2169 ^ n2162;
  assign n2327 = ~n2166 & n2326;
  assign n2328 = n2327 ^ n2169;
  assign n2321 = n2157 ^ n2061;
  assign n2322 = n2160 ^ n2061;
  assign n2323 = ~n2321 & n2322;
  assign n2324 = n2323 ^ n2157;
  assign n2316 = n2055 ^ n2052;
  assign n2317 = n2060 & ~n2316;
  assign n2318 = n2317 ^ n2052;
  assign n2309 = n2081 ^ n2068;
  assign n2310 = n2075 ^ n2068;
  assign n2311 = n2309 & ~n2310;
  assign n2312 = n2311 ^ n2081;
  assign n2304 = n2120 ^ n2113;
  assign n2305 = n2127 ^ n2113;
  assign n2306 = n2304 & ~n2305;
  assign n2307 = n2306 ^ n2120;
  assign n2301 = n2104 ^ n2090;
  assign n2302 = n2105 & ~n2301;
  assign n2303 = n2302 ^ n2097;
  assign n2308 = n2307 ^ n2303;
  assign n2313 = n2312 ^ n2308;
  assign n2298 = n2135 & ~n2142;
  assign n2290 = ~x14 & n618;
  assign n2291 = ~x13 & n622;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = x14 & n625;
  assign n2294 = x13 & n627;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = n2292 & n2295;
  assign n2283 = x22 & n166;
  assign n2284 = x21 & n168;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = ~x22 & n159;
  assign n2287 = ~x21 & n163;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = n2285 & n2288;
  assign n2297 = n2296 ^ n2289;
  assign n2299 = n2298 ^ n2297;
  assign n2273 = ~x16 & n460;
  assign n2274 = ~x15 & n462;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = x16 & n453;
  assign n2277 = x15 & n457;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n2275 & n2278;
  assign n2266 = ~x4 & n1734;
  assign n2267 = ~x3 & n1738;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = x4 & n1741;
  assign n2270 = x3 & n1743;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = n2268 & n2271;
  assign n2280 = n2279 ^ n2272;
  assign n2259 = ~x2 & n2013;
  assign n2260 = ~x1 & n2017;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = x2 & n2020;
  assign n2263 = x1 & n2022;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = n2261 & n2264;
  assign n2281 = n2280 ^ n2265;
  assign n2250 = x12 & n813;
  assign n2251 = x11 & n817;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = ~x12 & n820;
  assign n2254 = ~x11 & n822;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = n2252 & n2255;
  assign n2243 = x10 & n1044;
  assign n2244 = x9 & n1046;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = ~x10 & n1037;
  assign n2247 = ~x9 & n1041;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = n2245 & n2248;
  assign n2257 = n2256 ^ n2249;
  assign n2236 = ~x18 & n344;
  assign n2237 = ~x17 & n348;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = x18 & n351;
  assign n2240 = x17 & n353;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = n2238 & n2241;
  assign n2258 = n2257 ^ n2242;
  assign n2282 = n2281 ^ n2258;
  assign n2300 = n2299 ^ n2282;
  assign n2314 = n2313 ^ n2300;
  assign n2228 = ~x25 & n67;
  assign n2229 = n69 ^ x26;
  assign n2230 = n2229 ^ n69;
  assign n2231 = n71 & n2230;
  assign n2232 = n2231 ^ n69;
  assign n2233 = ~n2228 & ~n2232;
  assign n2220 = ~x8 & n1282;
  assign n2221 = ~x7 & n1284;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = x8 & n1275;
  assign n2224 = x7 & n1279;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = n2222 & n2225;
  assign n2213 = ~x6 & n1439;
  assign n2214 = ~x5 & n1443;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = x6 & n1446;
  assign n2217 = x5 & n1448;
  assign n2218 = ~n2216 & ~n2217;
  assign n2219 = n2215 & n2218;
  assign n2227 = n2226 ^ n2219;
  assign n2234 = n2233 ^ n2227;
  assign n2209 = n2032 ^ n2012;
  assign n2210 = n2033 & ~n2209;
  assign n2211 = n2210 ^ n2025;
  assign n2200 = ~x24 & n89;
  assign n2201 = ~x23 & n93;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = x24 & n96;
  assign n2204 = x23 & n98;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = n2202 & n2205;
  assign n2198 = x58 ^ x57;
  assign n2199 = x0 & n2198;
  assign n2207 = n2206 ^ n2199;
  assign n2191 = ~x20 & n225;
  assign n2192 = ~x19 & n229;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = x20 & n232;
  assign n2195 = x19 & n234;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = n2193 & n2196;
  assign n2208 = n2207 ^ n2197;
  assign n2212 = n2211 ^ n2208;
  assign n2235 = n2234 ^ n2212;
  assign n2315 = n2314 ^ n2235;
  assign n2319 = n2318 ^ n2315;
  assign n2187 = n2152 ^ n2131;
  assign n2188 = ~n2156 & n2187;
  assign n2189 = n2188 ^ n2131;
  assign n2182 = n2051 ^ n2043;
  assign n2183 = n2051 ^ n2046;
  assign n2184 = n2182 & n2183;
  assign n2185 = n2184 ^ n2043;
  assign n2178 = n2129 ^ n2083;
  assign n2179 = n2130 & ~n2178;
  assign n2180 = n2179 ^ n2106;
  assign n2174 = n2037 ^ n2034;
  assign n2175 = n2042 & ~n2174;
  assign n2176 = n2175 ^ n2034;
  assign n2171 = n2151 ^ n2147;
  assign n2172 = n2148 & ~n2171;
  assign n2173 = n2172 ^ n2143;
  assign n2177 = n2176 ^ n2173;
  assign n2181 = n2180 ^ n2177;
  assign n2186 = n2185 ^ n2181;
  assign n2190 = n2189 ^ n2186;
  assign n2320 = n2319 ^ n2190;
  assign n2325 = n2324 ^ n2320;
  assign n2329 = n2328 ^ n2325;
  assign n2502 = n2328 ^ n2320;
  assign n2503 = n2325 & n2502;
  assign n2504 = n2503 ^ n2328;
  assign n2497 = n2315 ^ n2190;
  assign n2498 = n2318 ^ n2190;
  assign n2499 = ~n2497 & n2498;
  assign n2500 = n2499 ^ n2315;
  assign n2492 = n2189 ^ n2185;
  assign n2493 = ~n2186 & n2492;
  assign n2494 = n2493 ^ n2181;
  assign n2487 = n2299 ^ n2281;
  assign n2488 = n2282 & n2487;
  assign n2489 = n2488 ^ n2258;
  assign n2476 = x23 & n166;
  assign n2477 = x22 & n168;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = ~x23 & n159;
  assign n2480 = ~x22 & n163;
  assign n2481 = ~n2479 & ~n2480;
  assign n2482 = n2478 & n2481;
  assign n2469 = x3 & n2020;
  assign n2470 = x2 & n2022;
  assign n2471 = ~n2469 & ~n2470;
  assign n2472 = ~x3 & n2013;
  assign n2473 = ~x2 & n2017;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = n2471 & n2474;
  assign n2483 = n2482 ^ n2475;
  assign n2456 = ~x59 & n2198;
  assign n2457 = x1 & n2456;
  assign n2458 = x59 ^ x58;
  assign n2459 = ~n2198 & n2458;
  assign n2460 = ~x59 & n2459;
  assign n2461 = x0 & n2460;
  assign n2462 = ~n2457 & ~n2461;
  assign n2463 = x59 & n2198;
  assign n2464 = ~x1 & n2463;
  assign n2465 = x59 & n2459;
  assign n2466 = ~x0 & n2465;
  assign n2467 = ~n2464 & ~n2466;
  assign n2468 = n2462 & n2467;
  assign n2484 = n2483 ^ n2468;
  assign n2447 = ~x13 & n820;
  assign n2448 = ~x12 & n822;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = x13 & n813;
  assign n2451 = x12 & n817;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = n2449 & n2452;
  assign n2440 = x21 & n232;
  assign n2441 = x20 & n234;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~x21 & n225;
  assign n2444 = ~x20 & n229;
  assign n2445 = ~n2443 & ~n2444;
  assign n2446 = n2442 & n2445;
  assign n2454 = n2453 ^ n2446;
  assign n2433 = ~x11 & n1037;
  assign n2434 = ~x10 & n1041;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = x11 & n1044;
  assign n2437 = x10 & n1046;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = n2435 & n2438;
  assign n2455 = n2454 ^ n2439;
  assign n2485 = n2484 ^ n2455;
  assign n2425 = ~x26 & n67;
  assign n2426 = n69 ^ x27;
  assign n2427 = n2426 ^ n69;
  assign n2428 = n71 & n2427;
  assign n2429 = n2428 ^ n69;
  assign n2430 = ~n2425 & ~n2429;
  assign n2418 = ~x17 & n460;
  assign n2419 = ~x16 & n462;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = x17 & n453;
  assign n2422 = x16 & n457;
  assign n2423 = ~n2421 & ~n2422;
  assign n2424 = n2420 & n2423;
  assign n2431 = n2430 ^ n2424;
  assign n2411 = ~x5 & n1734;
  assign n2412 = ~x4 & n1738;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = x5 & n1741;
  assign n2415 = x4 & n1743;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = n2413 & n2416;
  assign n2432 = n2431 ^ n2417;
  assign n2486 = n2485 ^ n2432;
  assign n2490 = n2489 ^ n2486;
  assign n2406 = n2298 ^ n2296;
  assign n2407 = n2297 & n2406;
  assign n2408 = n2407 ^ n2289;
  assign n2397 = ~x9 & n1282;
  assign n2398 = ~x8 & n1284;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = x9 & n1275;
  assign n2401 = x8 & n1279;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = n2399 & n2402;
  assign n2390 = x19 & n351;
  assign n2391 = x18 & n353;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~x19 & n344;
  assign n2394 = ~x18 & n348;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = n2392 & n2395;
  assign n2404 = n2403 ^ n2396;
  assign n2383 = ~x7 & n1439;
  assign n2384 = ~x6 & n1443;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = x7 & n1446;
  assign n2387 = x6 & n1448;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = n2385 & n2388;
  assign n2405 = n2404 ^ n2389;
  assign n2409 = n2408 ^ n2405;
  assign n2379 = n2206 ^ n2197;
  assign n2380 = ~n2207 & ~n2379;
  assign n2381 = n2380 ^ n2199;
  assign n2370 = ~x25 & n89;
  assign n2371 = ~x24 & n93;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = x25 & n96;
  assign n2374 = x24 & n98;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = n2372 & n2375;
  assign n2366 = x57 ^ x0;
  assign n2367 = ~n2198 & n2366;
  assign n2368 = n2367 ^ x0;
  assign n2369 = x59 & ~n2368;
  assign n2377 = n2376 ^ n2369;
  assign n2359 = x15 & n625;
  assign n2360 = x14 & n627;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~x15 & n618;
  assign n2363 = ~x14 & n622;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = n2361 & n2364;
  assign n2378 = n2377 ^ n2365;
  assign n2382 = n2381 ^ n2378;
  assign n2410 = n2409 ^ n2382;
  assign n2491 = n2490 ^ n2410;
  assign n2495 = n2494 ^ n2491;
  assign n2354 = n2180 ^ n2173;
  assign n2355 = ~n2177 & n2354;
  assign n2356 = n2355 ^ n2180;
  assign n2350 = n2300 ^ n2235;
  assign n2351 = n2313 ^ n2235;
  assign n2352 = n2350 & n2351;
  assign n2353 = n2352 ^ n2300;
  assign n2357 = n2356 ^ n2353;
  assign n2345 = n2312 ^ n2307;
  assign n2346 = n2308 & ~n2345;
  assign n2347 = n2346 ^ n2303;
  assign n2342 = n2234 ^ n2208;
  assign n2343 = n2212 & ~n2342;
  assign n2344 = n2343 ^ n2234;
  assign n2348 = n2347 ^ n2344;
  assign n2338 = n2279 ^ n2265;
  assign n2339 = n2280 & ~n2338;
  assign n2340 = n2339 ^ n2272;
  assign n2334 = n2233 ^ n2219;
  assign n2335 = ~n2227 & n2334;
  assign n2336 = n2335 ^ n2233;
  assign n2330 = n2249 ^ n2242;
  assign n2331 = n2256 ^ n2242;
  assign n2332 = n2330 & ~n2331;
  assign n2333 = n2332 ^ n2249;
  assign n2337 = n2336 ^ n2333;
  assign n2341 = n2340 ^ n2337;
  assign n2349 = n2348 ^ n2341;
  assign n2358 = n2357 ^ n2349;
  assign n2496 = n2495 ^ n2358;
  assign n2501 = n2500 ^ n2496;
  assign n2505 = n2504 ^ n2501;
  assign n2672 = n2504 ^ n2496;
  assign n2673 = ~n2501 & ~n2672;
  assign n2674 = n2673 ^ n2504;
  assign n2667 = n2491 ^ n2358;
  assign n2668 = n2494 ^ n2358;
  assign n2669 = n2667 & n2668;
  assign n2670 = n2669 ^ n2491;
  assign n2661 = n2353 ^ n2349;
  assign n2662 = n2356 ^ n2349;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n2663 ^ n2353;
  assign n2657 = n2344 ^ n2341;
  assign n2658 = ~n2348 & n2657;
  assign n2659 = n2658 ^ n2341;
  assign n2653 = n2408 ^ n2382;
  assign n2654 = n2409 & n2653;
  assign n2655 = n2654 ^ n2405;
  assign n2645 = ~x27 & n67;
  assign n2646 = n69 ^ x28;
  assign n2647 = n2646 ^ n69;
  assign n2648 = n71 & n2647;
  assign n2649 = n2648 ^ n69;
  assign n2650 = ~n2645 & ~n2649;
  assign n2637 = x8 & n1446;
  assign n2638 = x7 & n1448;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~x8 & n1439;
  assign n2641 = ~x7 & n1443;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = n2639 & n2642;
  assign n2630 = x10 & n1275;
  assign n2631 = x9 & n1279;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~x10 & n1282;
  assign n2634 = ~x9 & n1284;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = n2632 & n2635;
  assign n2644 = n2643 ^ n2636;
  assign n2651 = n2650 ^ n2644;
  assign n2620 = ~x2 & n2463;
  assign n2621 = ~x1 & n2465;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = x2 & n2456;
  assign n2624 = x1 & n2460;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = n2622 & n2625;
  assign n2613 = x24 & n166;
  assign n2614 = x23 & n168;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = ~x24 & n159;
  assign n2617 = ~x23 & n163;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = n2615 & n2618;
  assign n2627 = n2626 ^ n2619;
  assign n2606 = ~x16 & n618;
  assign n2607 = ~x15 & n622;
  assign n2608 = ~n2606 & ~n2607;
  assign n2609 = x16 & n625;
  assign n2610 = x15 & n627;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = n2608 & n2611;
  assign n2628 = n2627 ^ n2612;
  assign n2597 = ~x26 & n89;
  assign n2598 = ~x25 & n93;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = x26 & n96;
  assign n2601 = x25 & n98;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = n2599 & n2602;
  assign n2595 = x60 ^ x59;
  assign n2596 = x0 & n2595;
  assign n2604 = n2603 ^ n2596;
  assign n2588 = x22 & n232;
  assign n2589 = x21 & n234;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~x22 & n225;
  assign n2592 = ~x21 & n229;
  assign n2593 = ~n2591 & ~n2592;
  assign n2594 = n2590 & n2593;
  assign n2605 = n2604 ^ n2594;
  assign n2629 = n2628 ^ n2605;
  assign n2652 = n2651 ^ n2629;
  assign n2656 = n2655 ^ n2652;
  assign n2660 = n2659 ^ n2656;
  assign n2665 = n2664 ^ n2660;
  assign n2583 = n2486 ^ n2410;
  assign n2584 = n2489 ^ n2410;
  assign n2585 = ~n2583 & n2584;
  assign n2586 = n2585 ^ n2486;
  assign n2578 = n2381 ^ n2377;
  assign n2579 = n2378 & n2578;
  assign n2580 = n2579 ^ n2365;
  assign n2574 = n2340 ^ n2333;
  assign n2575 = ~n2337 & n2574;
  assign n2576 = n2575 ^ n2340;
  assign n2565 = ~x6 & n1734;
  assign n2566 = ~x5 & n1738;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = x6 & n1741;
  assign n2569 = x5 & n1743;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = n2567 & n2570;
  assign n2558 = x18 & n453;
  assign n2559 = x17 & n457;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~x18 & n460;
  assign n2562 = ~x17 & n462;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = n2560 & n2563;
  assign n2572 = n2571 ^ n2564;
  assign n2551 = ~x4 & n2013;
  assign n2552 = ~x3 & n2017;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = x4 & n2020;
  assign n2555 = x3 & n2022;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = n2553 & n2556;
  assign n2573 = n2572 ^ n2557;
  assign n2577 = n2576 ^ n2573;
  assign n2581 = n2580 ^ n2577;
  assign n2547 = n2455 ^ n2432;
  assign n2548 = ~n2485 & n2547;
  assign n2549 = n2548 ^ n2432;
  assign n2542 = n2403 ^ n2389;
  assign n2543 = n2404 & ~n2542;
  assign n2544 = n2543 ^ n2396;
  assign n2538 = n2453 ^ n2439;
  assign n2539 = n2454 & ~n2538;
  assign n2540 = n2539 ^ n2446;
  assign n2537 = n2369 & ~n2376;
  assign n2541 = n2540 ^ n2537;
  assign n2545 = n2544 ^ n2541;
  assign n2532 = n2482 ^ n2468;
  assign n2533 = n2483 & ~n2532;
  assign n2534 = n2533 ^ n2475;
  assign n2529 = n2424 ^ n2417;
  assign n2530 = n2431 & ~n2529;
  assign n2531 = n2530 ^ n2430;
  assign n2535 = n2534 ^ n2531;
  assign n2520 = ~x12 & n1037;
  assign n2521 = ~x11 & n1041;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = x12 & n1044;
  assign n2524 = x11 & n1046;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = n2522 & n2525;
  assign n2513 = ~x14 & n820;
  assign n2514 = ~x13 & n822;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = x14 & n813;
  assign n2517 = x13 & n817;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = n2515 & n2518;
  assign n2527 = n2526 ^ n2519;
  assign n2506 = ~x20 & n344;
  assign n2507 = ~x19 & n348;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = x20 & n351;
  assign n2510 = x19 & n353;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = n2508 & n2511;
  assign n2528 = n2527 ^ n2512;
  assign n2536 = n2535 ^ n2528;
  assign n2546 = n2545 ^ n2536;
  assign n2550 = n2549 ^ n2546;
  assign n2582 = n2581 ^ n2550;
  assign n2587 = n2586 ^ n2582;
  assign n2666 = n2665 ^ n2587;
  assign n2671 = n2670 ^ n2666;
  assign n2675 = n2674 ^ n2671;
  assign n2860 = n2674 ^ n2666;
  assign n2861 = ~n2671 & n2860;
  assign n2862 = n2861 ^ n2674;
  assign n2856 = n2660 ^ n2587;
  assign n2857 = ~n2665 & n2856;
  assign n2858 = n2857 ^ n2587;
  assign n2851 = n2659 ^ n2655;
  assign n2852 = ~n2656 & ~n2851;
  assign n2853 = n2852 ^ n2652;
  assign n2848 = n2586 ^ n2581;
  assign n2849 = ~n2582 & ~n2848;
  assign n2850 = n2849 ^ n2550;
  assign n2854 = n2853 ^ n2850;
  assign n2843 = n2549 ^ n2536;
  assign n2844 = n2546 & n2843;
  assign n2845 = n2844 ^ n2549;
  assign n2838 = n2580 ^ n2573;
  assign n2839 = n2580 ^ n2576;
  assign n2840 = n2838 & ~n2839;
  assign n2841 = n2840 ^ n2573;
  assign n2827 = ~x21 & n344;
  assign n2828 = ~x20 & n348;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = x21 & n351;
  assign n2831 = x20 & n353;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = n2829 & n2832;
  assign n2820 = ~x13 & n1037;
  assign n2821 = ~x12 & n1041;
  assign n2822 = ~n2820 & ~n2821;
  assign n2823 = x13 & n1044;
  assign n2824 = x12 & n1046;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = n2822 & n2825;
  assign n2834 = n2833 ^ n2826;
  assign n2813 = x11 & n1275;
  assign n2814 = x10 & n1279;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = ~x11 & n1282;
  assign n2817 = ~x10 & n1284;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = n2815 & n2818;
  assign n2835 = n2834 ^ n2819;
  assign n2804 = ~x5 & n2013;
  assign n2805 = ~x4 & n2017;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = x5 & n2020;
  assign n2808 = x4 & n2022;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = n2806 & n2809;
  assign n2797 = ~x7 & n1734;
  assign n2798 = ~x6 & n1738;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = x7 & n1741;
  assign n2801 = x6 & n1743;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n2799 & n2802;
  assign n2811 = n2810 ^ n2803;
  assign n2790 = ~x17 & n618;
  assign n2791 = ~x16 & n622;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = x17 & n625;
  assign n2794 = x16 & n627;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = n2792 & n2795;
  assign n2812 = n2811 ^ n2796;
  assign n2836 = n2835 ^ n2812;
  assign n2781 = x25 & n166;
  assign n2782 = x24 & n168;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~x25 & n159;
  assign n2785 = ~x24 & n163;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = n2783 & n2786;
  assign n2774 = ~x9 & n1439;
  assign n2775 = ~x8 & n1443;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = x9 & n1446;
  assign n2778 = x8 & n1448;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = n2776 & n2779;
  assign n2788 = n2787 ^ n2780;
  assign n2767 = ~x19 & n460;
  assign n2768 = ~x18 & n462;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = x19 & n453;
  assign n2771 = x18 & n457;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = n2769 & n2772;
  assign n2789 = n2788 ^ n2773;
  assign n2837 = n2836 ^ n2789;
  assign n2842 = n2841 ^ n2837;
  assign n2846 = n2845 ^ n2842;
  assign n2761 = n2651 ^ n2605;
  assign n2762 = n2651 ^ n2628;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = n2763 ^ n2605;
  assign n2757 = n2544 ^ n2540;
  assign n2758 = ~n2541 & ~n2757;
  assign n2759 = n2758 ^ n2537;
  assign n2742 = x61 & n2595;
  assign n2743 = ~x1 & n2742;
  assign n2744 = x61 ^ x60;
  assign n2745 = ~n2595 & n2744;
  assign n2746 = x61 & n2745;
  assign n2747 = ~x0 & n2746;
  assign n2748 = ~n2743 & ~n2747;
  assign n2749 = ~x61 & n2595;
  assign n2750 = x1 & n2749;
  assign n2751 = ~x61 & n2745;
  assign n2752 = x0 & n2751;
  assign n2753 = ~n2750 & ~n2752;
  assign n2754 = n2748 & n2753;
  assign n2735 = x3 & n2456;
  assign n2736 = x2 & n2460;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = ~x3 & n2463;
  assign n2739 = ~x2 & n2465;
  assign n2740 = ~n2738 & ~n2739;
  assign n2741 = n2737 & n2740;
  assign n2755 = n2754 ^ n2741;
  assign n2728 = ~x28 & n67;
  assign n2729 = n69 ^ x29;
  assign n2730 = n2729 ^ n69;
  assign n2731 = n71 & n2730;
  assign n2732 = n2731 ^ n69;
  assign n2733 = ~n2728 & ~n2732;
  assign n2724 = x59 ^ x0;
  assign n2725 = ~n2595 & n2724;
  assign n2726 = n2725 ^ x0;
  assign n2727 = x61 & ~n2726;
  assign n2734 = n2733 ^ n2727;
  assign n2756 = n2755 ^ n2734;
  assign n2760 = n2759 ^ n2756;
  assign n2765 = n2764 ^ n2760;
  assign n2719 = n2531 ^ n2528;
  assign n2720 = ~n2535 & n2719;
  assign n2721 = n2720 ^ n2528;
  assign n2715 = n2526 ^ n2512;
  assign n2716 = n2527 & ~n2715;
  assign n2717 = n2716 ^ n2519;
  assign n2711 = n2650 ^ n2636;
  assign n2712 = ~n2644 & n2711;
  assign n2713 = n2712 ^ n2650;
  assign n2707 = n2596 ^ n2594;
  assign n2708 = n2603 ^ n2594;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = n2709 ^ n2596;
  assign n2714 = n2713 ^ n2710;
  assign n2718 = n2717 ^ n2714;
  assign n2722 = n2721 ^ n2718;
  assign n2702 = n2619 ^ n2612;
  assign n2703 = ~n2627 & n2702;
  assign n2704 = n2703 ^ n2612;
  assign n2699 = n2564 ^ n2557;
  assign n2700 = ~n2572 & n2699;
  assign n2701 = n2700 ^ n2557;
  assign n2705 = n2704 ^ n2701;
  assign n2690 = ~x23 & n225;
  assign n2691 = ~x22 & n229;
  assign n2692 = ~n2690 & ~n2691;
  assign n2693 = x23 & n232;
  assign n2694 = x22 & n234;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = n2692 & n2695;
  assign n2683 = x27 & n96;
  assign n2684 = x26 & n98;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~x27 & n89;
  assign n2687 = ~x26 & n93;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = n2685 & n2688;
  assign n2697 = n2696 ^ n2689;
  assign n2676 = ~x15 & n820;
  assign n2677 = ~x14 & n822;
  assign n2678 = ~n2676 & ~n2677;
  assign n2679 = x15 & n813;
  assign n2680 = x14 & n817;
  assign n2681 = ~n2679 & ~n2680;
  assign n2682 = n2678 & n2681;
  assign n2698 = n2697 ^ n2682;
  assign n2706 = n2705 ^ n2698;
  assign n2723 = n2722 ^ n2706;
  assign n2766 = n2765 ^ n2723;
  assign n2847 = n2846 ^ n2766;
  assign n2855 = n2854 ^ n2847;
  assign n2859 = n2858 ^ n2855;
  assign n2863 = n2862 ^ n2859;
  assign n3041 = n2862 ^ n2855;
  assign n3042 = ~n2859 & n3041;
  assign n3043 = n3042 ^ n2862;
  assign n3037 = n2850 ^ n2847;
  assign n3038 = ~n2854 & n3037;
  assign n3039 = n3038 ^ n2847;
  assign n3033 = n2846 ^ n2765;
  assign n3034 = ~n2766 & ~n3033;
  assign n3035 = n3034 ^ n2723;
  assign n3027 = n2845 ^ n2837;
  assign n3028 = n2845 ^ n2841;
  assign n3029 = n3027 & ~n3028;
  assign n3030 = n3029 ^ n2837;
  assign n3022 = n2812 ^ n2789;
  assign n3023 = ~n2836 & n3022;
  assign n3024 = n3023 ^ n2789;
  assign n3018 = n2717 ^ n2710;
  assign n3019 = n2714 & ~n3018;
  assign n3020 = n3019 ^ n2717;
  assign n3014 = n2696 ^ n2682;
  assign n3015 = n2697 & ~n3014;
  assign n3016 = n3015 ^ n2689;
  assign n3012 = n2727 & ~n2733;
  assign n3005 = ~x2 & n2742;
  assign n3006 = ~x1 & n2746;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = x2 & n2749;
  assign n3009 = x1 & n2751;
  assign n3010 = ~n3008 & ~n3009;
  assign n3011 = n3007 & n3010;
  assign n3013 = n3012 ^ n3011;
  assign n3017 = n3016 ^ n3013;
  assign n3021 = n3020 ^ n3017;
  assign n3025 = n3024 ^ n3021;
  assign n3000 = n2701 ^ n2698;
  assign n3001 = ~n2705 & n3000;
  assign n3002 = n3001 ^ n2698;
  assign n2996 = n2810 ^ n2796;
  assign n2997 = n2811 & ~n2996;
  assign n2998 = n2997 ^ n2803;
  assign n2992 = n2833 ^ n2819;
  assign n2993 = n2834 & ~n2992;
  assign n2994 = n2993 ^ n2826;
  assign n2989 = n2787 ^ n2773;
  assign n2990 = n2788 & ~n2989;
  assign n2991 = n2990 ^ n2780;
  assign n2995 = n2994 ^ n2991;
  assign n2999 = n2998 ^ n2995;
  assign n3003 = n3002 ^ n2999;
  assign n2985 = n2754 ^ n2734;
  assign n2986 = n2755 & ~n2985;
  assign n2987 = n2986 ^ n2741;
  assign n2975 = ~x12 & n1282;
  assign n2976 = ~x11 & n1284;
  assign n2977 = ~n2975 & ~n2976;
  assign n2978 = x12 & n1275;
  assign n2979 = x11 & n1279;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n2977 & n2980;
  assign n2968 = ~x22 & n344;
  assign n2969 = ~x21 & n348;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = x22 & n351;
  assign n2972 = x21 & n353;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = n2970 & n2973;
  assign n2982 = n2981 ^ n2974;
  assign n2961 = ~x10 & n1439;
  assign n2962 = ~x9 & n1443;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = x10 & n1446;
  assign n2965 = x9 & n1448;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = n2963 & n2966;
  assign n2983 = n2982 ^ n2967;
  assign n2952 = ~x16 & n820;
  assign n2953 = ~x15 & n822;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = x16 & n813;
  assign n2956 = x15 & n817;
  assign n2957 = ~n2955 & ~n2956;
  assign n2958 = n2954 & n2957;
  assign n2945 = x24 & n232;
  assign n2946 = x23 & n234;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~x24 & n225;
  assign n2949 = ~x23 & n229;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n2947 & n2950;
  assign n2959 = n2958 ^ n2951;
  assign n2938 = ~x14 & n1037;
  assign n2939 = ~x13 & n1041;
  assign n2940 = ~n2938 & ~n2939;
  assign n2941 = x14 & n1044;
  assign n2942 = x13 & n1046;
  assign n2943 = ~n2941 & ~n2942;
  assign n2944 = n2940 & n2943;
  assign n2960 = n2959 ^ n2944;
  assign n2984 = n2983 ^ n2960;
  assign n2988 = n2987 ^ n2984;
  assign n3004 = n3003 ^ n2988;
  assign n3026 = n3025 ^ n3004;
  assign n3031 = n3030 ^ n3026;
  assign n2933 = n2764 ^ n2756;
  assign n2934 = n2764 ^ n2759;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n2935 ^ n2756;
  assign n2929 = n2718 ^ n2706;
  assign n2930 = n2722 & ~n2929;
  assign n2931 = n2930 ^ n2706;
  assign n2918 = ~x18 & n618;
  assign n2919 = ~x17 & n622;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = x18 & n625;
  assign n2922 = x17 & n627;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = n2920 & n2923;
  assign n2911 = ~x6 & n2013;
  assign n2912 = ~x5 & n2017;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = x6 & n2020;
  assign n2915 = x5 & n2022;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = n2913 & n2916;
  assign n2925 = n2924 ^ n2917;
  assign n2904 = x4 & n2456;
  assign n2905 = x3 & n2460;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = ~x4 & n2463;
  assign n2908 = ~x3 & n2465;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = n2906 & n2909;
  assign n2926 = n2925 ^ n2910;
  assign n2896 = ~x28 & n89;
  assign n2897 = ~x27 & n93;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = x28 & n96;
  assign n2900 = x27 & n98;
  assign n2901 = ~n2899 & ~n2900;
  assign n2902 = n2898 & n2901;
  assign n2889 = ~x29 & n67;
  assign n2890 = n69 ^ x30;
  assign n2891 = n2890 ^ n69;
  assign n2892 = n71 & n2891;
  assign n2893 = n2892 ^ n69;
  assign n2894 = ~n2889 & ~n2893;
  assign n2887 = x62 ^ x61;
  assign n2888 = x0 & n2887;
  assign n2895 = n2894 ^ n2888;
  assign n2903 = n2902 ^ n2895;
  assign n2927 = n2926 ^ n2903;
  assign n2878 = ~x20 & n460;
  assign n2879 = ~x19 & n462;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = x20 & n453;
  assign n2882 = x19 & n457;
  assign n2883 = ~n2881 & ~n2882;
  assign n2884 = n2880 & n2883;
  assign n2871 = ~x26 & n159;
  assign n2872 = ~x25 & n163;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = x26 & n166;
  assign n2875 = x25 & n168;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = n2873 & n2876;
  assign n2885 = n2884 ^ n2877;
  assign n2864 = x8 & n1741;
  assign n2865 = x7 & n1743;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = ~x8 & n1734;
  assign n2868 = ~x7 & n1738;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = n2866 & n2869;
  assign n2886 = n2885 ^ n2870;
  assign n2928 = n2927 ^ n2886;
  assign n2932 = n2931 ^ n2928;
  assign n2937 = n2936 ^ n2932;
  assign n3032 = n3031 ^ n2937;
  assign n3036 = n3035 ^ n3032;
  assign n3040 = n3039 ^ n3036;
  assign n3044 = n3043 ^ n3040;
  assign n3241 = n3043 ^ n3036;
  assign n3242 = ~n3040 & n3241;
  assign n3243 = n3242 ^ n3043;
  assign n3236 = n3035 ^ n2937;
  assign n3237 = n3035 ^ n3031;
  assign n3238 = n3236 & ~n3237;
  assign n3239 = n3238 ^ n2937;
  assign n3232 = n3030 ^ n3025;
  assign n3233 = ~n3026 & n3232;
  assign n3234 = n3233 ^ n3004;
  assign n3227 = n2936 ^ n2931;
  assign n3228 = ~n2932 & ~n3227;
  assign n3229 = n3228 ^ n2928;
  assign n3221 = n2987 ^ n2983;
  assign n3222 = n2984 & ~n3221;
  assign n3223 = n3222 ^ n2960;
  assign n3217 = n2903 ^ n2886;
  assign n3218 = n2926 ^ n2886;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = n3219 ^ n2903;
  assign n3224 = n3223 ^ n3220;
  assign n3206 = x19 & n625;
  assign n3207 = x18 & n627;
  assign n3208 = ~n3206 & ~n3207;
  assign n3209 = ~x19 & n618;
  assign n3210 = ~x18 & n622;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = n3208 & n3211;
  assign n3199 = ~x5 & n2463;
  assign n3200 = ~x4 & n2465;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = x5 & n2456;
  assign n3203 = x4 & n2460;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = n3201 & n3204;
  assign n3213 = n3212 ^ n3205;
  assign n3192 = ~x3 & n2742;
  assign n3193 = ~x2 & n2746;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = x3 & n2749;
  assign n3196 = x2 & n2751;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = n3194 & n3197;
  assign n3214 = n3213 ^ n3198;
  assign n3183 = ~x25 & n225;
  assign n3184 = ~x24 & n229;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = x25 & n232;
  assign n3187 = x24 & n234;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = n3185 & n3188;
  assign n3176 = ~x29 & n89;
  assign n3177 = ~x28 & n93;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = x29 & n96;
  assign n3180 = x28 & n98;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = n3178 & n3181;
  assign n3190 = n3189 ^ n3182;
  assign n3163 = x63 & n2887;
  assign n3164 = ~x1 & n3163;
  assign n3165 = x63 ^ x62;
  assign n3166 = ~n2887 & n3165;
  assign n3167 = x63 & n3166;
  assign n3168 = ~x0 & n3167;
  assign n3169 = ~n3164 & ~n3168;
  assign n3170 = ~x63 & n2887;
  assign n3171 = x1 & n3170;
  assign n3172 = ~x63 & n3166;
  assign n3173 = x0 & n3172;
  assign n3174 = ~n3171 & ~n3173;
  assign n3175 = n3169 & n3174;
  assign n3191 = n3190 ^ n3175;
  assign n3215 = n3214 ^ n3191;
  assign n3154 = x17 & n813;
  assign n3155 = x16 & n817;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = ~x17 & n820;
  assign n3158 = ~x16 & n822;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = n3156 & n3159;
  assign n3147 = ~x15 & n1037;
  assign n3148 = ~x14 & n1041;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = x15 & n1044;
  assign n3151 = x14 & n1046;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = n3149 & n3152;
  assign n3161 = n3160 ^ n3153;
  assign n3140 = ~x23 & n344;
  assign n3141 = ~x22 & n348;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = x23 & n351;
  assign n3144 = x22 & n353;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = n3142 & n3145;
  assign n3162 = n3161 ^ n3146;
  assign n3216 = n3215 ^ n3162;
  assign n3225 = n3224 ^ n3216;
  assign n3135 = n3016 ^ n3012;
  assign n3136 = ~n3013 & n3135;
  assign n3137 = n3136 ^ n3011;
  assign n3131 = n2924 ^ n2910;
  assign n3132 = n2925 & ~n3131;
  assign n3133 = n3132 ^ n2917;
  assign n3127 = n2884 ^ n2870;
  assign n3128 = n2885 & ~n3127;
  assign n3129 = n3128 ^ n2877;
  assign n3124 = n2981 ^ n2967;
  assign n3125 = n2982 & ~n3124;
  assign n3126 = n3125 ^ n2974;
  assign n3130 = n3129 ^ n3126;
  assign n3134 = n3133 ^ n3130;
  assign n3138 = n3137 ^ n3134;
  assign n3120 = n2958 ^ n2944;
  assign n3121 = n2959 & ~n3120;
  assign n3122 = n3121 ^ n2951;
  assign n3116 = n2902 ^ n2894;
  assign n3117 = ~n2895 & ~n3116;
  assign n3118 = n3117 ^ n2888;
  assign n3109 = ~x30 & n67;
  assign n3110 = n69 ^ x31;
  assign n3111 = n3110 ^ n69;
  assign n3112 = n71 & n3111;
  assign n3113 = n3112 ^ n69;
  assign n3114 = ~n3109 & ~n3113;
  assign n3105 = x61 ^ x0;
  assign n3106 = ~n2887 & n3105;
  assign n3107 = n3106 ^ x0;
  assign n3108 = x63 & ~n3107;
  assign n3115 = n3114 ^ n3108;
  assign n3119 = n3118 ^ n3115;
  assign n3123 = n3122 ^ n3119;
  assign n3139 = n3138 ^ n3123;
  assign n3226 = n3225 ^ n3139;
  assign n3230 = n3229 ^ n3226;
  assign n3101 = n2999 ^ n2988;
  assign n3102 = ~n3003 & n3101;
  assign n3103 = n3102 ^ n2988;
  assign n3096 = n3024 ^ n3017;
  assign n3097 = n3024 ^ n3020;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n3098 ^ n3017;
  assign n3092 = n2998 ^ n2991;
  assign n3093 = ~n2995 & n3092;
  assign n3094 = n3093 ^ n2998;
  assign n3082 = ~x11 & n1439;
  assign n3083 = ~x10 & n1443;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = x11 & n1446;
  assign n3086 = x10 & n1448;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = n3084 & n3087;
  assign n3075 = x13 & n1275;
  assign n3076 = x12 & n1279;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~x13 & n1282;
  assign n3079 = ~x12 & n1284;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = n3077 & n3080;
  assign n3089 = n3088 ^ n3081;
  assign n3068 = ~x27 & n159;
  assign n3069 = ~x26 & n163;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = x27 & n166;
  assign n3072 = x26 & n168;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = n3070 & n3073;
  assign n3090 = n3089 ^ n3074;
  assign n3059 = x21 & n453;
  assign n3060 = x20 & n457;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = ~x21 & n460;
  assign n3063 = ~x20 & n462;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n3061 & n3064;
  assign n3052 = ~x9 & n1734;
  assign n3053 = ~x8 & n1738;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = x9 & n1741;
  assign n3056 = x8 & n1743;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = n3054 & n3057;
  assign n3066 = n3065 ^ n3058;
  assign n3045 = x7 & n2020;
  assign n3046 = x6 & n2022;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = ~x7 & n2013;
  assign n3049 = ~x6 & n2017;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = n3047 & n3050;
  assign n3067 = n3066 ^ n3051;
  assign n3091 = n3090 ^ n3067;
  assign n3095 = n3094 ^ n3091;
  assign n3100 = n3099 ^ n3095;
  assign n3104 = n3103 ^ n3100;
  assign n3231 = n3230 ^ n3104;
  assign n3235 = n3234 ^ n3231;
  assign n3240 = n3239 ^ n3235;
  assign n3244 = n3243 ^ n3240;
  assign n3428 = n3243 ^ n3235;
  assign n3429 = n3240 & ~n3428;
  assign n3430 = n3429 ^ n3243;
  assign n3424 = n3234 ^ n3230;
  assign n3425 = n3231 & n3424;
  assign n3426 = n3425 ^ n3104;
  assign n3419 = n3229 ^ n3225;
  assign n3420 = n3226 & ~n3419;
  assign n3421 = n3420 ^ n3139;
  assign n3416 = n3103 ^ n3099;
  assign n3417 = ~n3100 & n3416;
  assign n3418 = n3417 ^ n3095;
  assign n3422 = n3421 ^ n3418;
  assign n3411 = n3220 ^ n3216;
  assign n3412 = n3224 & ~n3411;
  assign n3413 = n3412 ^ n3216;
  assign n3407 = n3134 ^ n3123;
  assign n3408 = ~n3138 & ~n3407;
  assign n3409 = n3408 ^ n3123;
  assign n3403 = n3133 ^ n3129;
  assign n3404 = n3130 & ~n3403;
  assign n3405 = n3404 ^ n3126;
  assign n3393 = ~x26 & n225;
  assign n3394 = ~x25 & n229;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = x26 & n232;
  assign n3397 = x25 & n234;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = n3395 & n3398;
  assign n3386 = x2 & n3170;
  assign n3387 = x1 & n3172;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = ~x2 & n3163;
  assign n3390 = ~x1 & n3167;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = n3388 & n3391;
  assign n3400 = n3399 ^ n3392;
  assign n3379 = x18 & n813;
  assign n3380 = x17 & n817;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = ~x18 & n820;
  assign n3383 = ~x17 & n822;
  assign n3384 = ~n3382 & ~n3383;
  assign n3385 = n3381 & n3384;
  assign n3401 = n3400 ^ n3385;
  assign n3370 = ~x4 & n2742;
  assign n3371 = ~x3 & n2746;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = x4 & n2749;
  assign n3374 = x3 & n2751;
  assign n3375 = ~n3373 & ~n3374;
  assign n3376 = n3372 & n3375;
  assign n3363 = ~x6 & n2463;
  assign n3364 = ~x5 & n2465;
  assign n3365 = ~n3363 & ~n3364;
  assign n3366 = x6 & n2456;
  assign n3367 = x5 & n2460;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = n3365 & n3368;
  assign n3377 = n3376 ^ n3369;
  assign n3362 = n3108 & ~n3114;
  assign n3378 = n3377 ^ n3362;
  assign n3402 = n3401 ^ n3378;
  assign n3406 = n3405 ^ n3402;
  assign n3410 = n3409 ^ n3406;
  assign n3414 = n3413 ^ n3410;
  assign n3357 = n3094 ^ n3090;
  assign n3358 = n3091 & ~n3357;
  assign n3359 = n3358 ^ n3067;
  assign n3351 = n3081 ^ n3074;
  assign n3352 = n3088 ^ n3074;
  assign n3353 = n3351 & ~n3352;
  assign n3354 = n3353 ^ n3081;
  assign n3347 = n3189 ^ n3175;
  assign n3348 = n3190 & ~n3347;
  assign n3349 = n3348 ^ n3182;
  assign n3344 = n3153 ^ n3146;
  assign n3345 = ~n3161 & n3344;
  assign n3346 = n3345 ^ n3146;
  assign n3350 = n3349 ^ n3346;
  assign n3355 = n3354 ^ n3350;
  assign n3333 = x12 & n1446;
  assign n3334 = x11 & n1448;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~x12 & n1439;
  assign n3337 = ~x11 & n1443;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = n3335 & n3338;
  assign n3326 = x28 & n166;
  assign n3327 = x27 & n168;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~x28 & n159;
  assign n3330 = ~x27 & n163;
  assign n3331 = ~n3329 & ~n3330;
  assign n3332 = n3328 & n3331;
  assign n3340 = n3339 ^ n3332;
  assign n3319 = x22 & n453;
  assign n3320 = x21 & n457;
  assign n3321 = ~n3319 & ~n3320;
  assign n3322 = ~x22 & n460;
  assign n3323 = ~x21 & n462;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = n3321 & n3324;
  assign n3341 = n3340 ^ n3325;
  assign n3310 = ~x16 & n1037;
  assign n3311 = ~x15 & n1041;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = x16 & n1044;
  assign n3314 = x15 & n1046;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = n3312 & n3315;
  assign n3303 = ~x24 & n344;
  assign n3304 = ~x23 & n348;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = x24 & n351;
  assign n3307 = x23 & n353;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = n3305 & n3308;
  assign n3317 = n3316 ^ n3309;
  assign n3296 = ~x14 & n1282;
  assign n3297 = ~x13 & n1284;
  assign n3298 = ~n3296 & ~n3297;
  assign n3299 = x14 & n1275;
  assign n3300 = x13 & n1279;
  assign n3301 = ~n3299 & ~n3300;
  assign n3302 = n3298 & n3301;
  assign n3318 = n3317 ^ n3302;
  assign n3342 = n3341 ^ n3318;
  assign n3287 = x8 & n2020;
  assign n3288 = x7 & n2022;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = ~x8 & n2013;
  assign n3291 = ~x7 & n2017;
  assign n3292 = ~n3290 & ~n3291;
  assign n3293 = n3289 & n3292;
  assign n3280 = ~x10 & n1734;
  assign n3281 = ~x9 & n1738;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = x10 & n1741;
  assign n3284 = x9 & n1743;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286 = n3282 & n3285;
  assign n3294 = n3293 ^ n3286;
  assign n3273 = x20 & n625;
  assign n3274 = x19 & n627;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = ~x20 & n618;
  assign n3277 = ~x19 & n622;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = n3275 & n3278;
  assign n3295 = n3294 ^ n3279;
  assign n3343 = n3342 ^ n3295;
  assign n3356 = n3355 ^ n3343;
  assign n3360 = n3359 ^ n3356;
  assign n3268 = n3122 ^ n3118;
  assign n3269 = ~n3119 & n3268;
  assign n3270 = n3269 ^ n3115;
  assign n3265 = n3191 ^ n3162;
  assign n3266 = ~n3215 & n3265;
  assign n3267 = n3266 ^ n3162;
  assign n3271 = n3270 ^ n3267;
  assign n3260 = n3205 ^ n3198;
  assign n3261 = ~n3213 & n3260;
  assign n3262 = n3261 ^ n3198;
  assign n3257 = n3058 ^ n3051;
  assign n3258 = ~n3066 & n3257;
  assign n3259 = n3258 ^ n3051;
  assign n3263 = n3262 ^ n3259;
  assign n3249 = ~x30 & n89;
  assign n3250 = ~x29 & n93;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = x30 & n96;
  assign n3253 = x29 & n98;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = n3251 & n3254;
  assign n3246 = x31 & n67;
  assign n3247 = n3246 ^ x33;
  assign n3245 = x0 & x63;
  assign n3248 = n3247 ^ n3245;
  assign n3256 = n3255 ^ n3248;
  assign n3264 = n3263 ^ n3256;
  assign n3272 = n3271 ^ n3264;
  assign n3361 = n3360 ^ n3272;
  assign n3415 = n3414 ^ n3361;
  assign n3423 = n3422 ^ n3415;
  assign n3427 = n3426 ^ n3423;
  assign n3431 = n3430 ^ n3427;
  assign n3618 = n3430 ^ n3423;
  assign n3619 = ~n3427 & n3618;
  assign n3620 = n3619 ^ n3430;
  assign n3614 = n3418 ^ n3415;
  assign n3615 = n3422 & n3614;
  assign n3616 = n3615 ^ n3415;
  assign n3610 = n3414 ^ n3360;
  assign n3611 = n3361 & ~n3610;
  assign n3612 = n3611 ^ n3272;
  assign n3605 = n3413 ^ n3409;
  assign n3606 = n3410 & n3605;
  assign n3607 = n3606 ^ n3406;
  assign n3601 = n3359 ^ n3355;
  assign n3602 = n3356 & ~n3601;
  assign n3603 = n3602 ^ n3343;
  assign n3597 = n3405 ^ n3401;
  assign n3598 = ~n3402 & ~n3597;
  assign n3599 = n3598 ^ n3378;
  assign n3590 = n3332 ^ n3325;
  assign n3591 = n3339 ^ n3325;
  assign n3592 = n3590 & ~n3591;
  assign n3593 = n3592 ^ n3332;
  assign n3581 = ~x3 & n3163;
  assign n3582 = ~x2 & n3167;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = x3 & n3170;
  assign n3585 = x2 & n3172;
  assign n3586 = ~n3584 & ~n3585;
  assign n3587 = n3583 & n3586;
  assign n3574 = ~x19 & n820;
  assign n3575 = ~x18 & n822;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = x19 & n813;
  assign n3578 = x18 & n817;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = n3576 & n3579;
  assign n3588 = n3587 ^ n3580;
  assign n3573 = x1 & x63;
  assign n3589 = n3588 ^ n3573;
  assign n3594 = n3593 ^ n3589;
  assign n3564 = ~x9 & n2013;
  assign n3565 = ~x8 & n2017;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = x9 & n2020;
  assign n3568 = x8 & n2022;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = n3566 & n3569;
  assign n3557 = ~x21 & n618;
  assign n3558 = ~x20 & n622;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = x21 & n625;
  assign n3561 = x20 & n627;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = n3559 & n3562;
  assign n3571 = n3570 ^ n3563;
  assign n3550 = x7 & n2456;
  assign n3551 = x6 & n2460;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = ~x7 & n2463;
  assign n3554 = ~x6 & n2465;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = n3552 & n3555;
  assign n3572 = n3571 ^ n3556;
  assign n3595 = n3594 ^ n3572;
  assign n3539 = ~x17 & n1037;
  assign n3540 = ~x16 & n1041;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = x17 & n1044;
  assign n3543 = x16 & n1046;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = n3541 & n3544;
  assign n3532 = ~x31 & n89;
  assign n3533 = ~x30 & n93;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = x31 & n96;
  assign n3536 = x30 & n98;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = n3534 & n3537;
  assign n3546 = n3545 ^ n3538;
  assign n3525 = x27 & n232;
  assign n3526 = x26 & n234;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = ~x27 & n225;
  assign n3529 = ~x26 & n229;
  assign n3530 = ~n3528 & ~n3529;
  assign n3531 = n3527 & n3530;
  assign n3547 = n3546 ^ n3531;
  assign n3516 = x23 & n453;
  assign n3517 = x22 & n457;
  assign n3518 = ~n3516 & ~n3517;
  assign n3519 = ~x23 & n460;
  assign n3520 = ~x22 & n462;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = n3518 & n3521;
  assign n3509 = ~x29 & n159;
  assign n3510 = ~x28 & n163;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = x29 & n166;
  assign n3513 = x28 & n168;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = n3511 & n3514;
  assign n3523 = n3522 ^ n3515;
  assign n3502 = ~x11 & n1734;
  assign n3503 = ~x10 & n1738;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = x11 & n1741;
  assign n3506 = x10 & n1743;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = n3504 & n3507;
  assign n3524 = n3523 ^ n3508;
  assign n3548 = n3547 ^ n3524;
  assign n3493 = ~x25 & n344;
  assign n3494 = ~x24 & n348;
  assign n3495 = ~n3493 & ~n3494;
  assign n3496 = x25 & n351;
  assign n3497 = x24 & n353;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = n3495 & n3498;
  assign n3486 = x15 & n1275;
  assign n3487 = x14 & n1279;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = ~x15 & n1282;
  assign n3490 = ~x14 & n1284;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = n3488 & n3491;
  assign n3500 = n3499 ^ n3492;
  assign n3479 = ~x13 & n1439;
  assign n3480 = ~x12 & n1443;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = x13 & n1446;
  assign n3483 = x12 & n1448;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = n3481 & n3484;
  assign n3501 = n3500 ^ n3485;
  assign n3549 = n3548 ^ n3501;
  assign n3596 = n3595 ^ n3549;
  assign n3600 = n3599 ^ n3596;
  assign n3604 = n3603 ^ n3600;
  assign n3608 = n3607 ^ n3604;
  assign n3473 = n3267 ^ n3264;
  assign n3474 = n3270 ^ n3264;
  assign n3475 = n3473 & ~n3474;
  assign n3476 = n3475 ^ n3267;
  assign n3469 = n3259 ^ n3256;
  assign n3470 = ~n3263 & n3469;
  assign n3471 = n3470 ^ n3256;
  assign n3465 = n3354 ^ n3349;
  assign n3466 = n3350 & ~n3465;
  assign n3467 = n3466 ^ n3346;
  assign n3462 = n3376 ^ n3362;
  assign n3463 = n3377 & n3462;
  assign n3464 = n3463 ^ n3369;
  assign n3468 = n3467 ^ n3464;
  assign n3472 = n3471 ^ n3468;
  assign n3477 = n3476 ^ n3472;
  assign n3458 = n3341 ^ n3295;
  assign n3459 = n3342 & ~n3458;
  assign n3460 = n3459 ^ n3318;
  assign n3452 = n3286 ^ n3279;
  assign n3453 = n3293 ^ n3279;
  assign n3454 = n3452 & ~n3453;
  assign n3455 = n3454 ^ n3286;
  assign n3448 = n3316 ^ n3302;
  assign n3449 = n3317 & ~n3448;
  assign n3450 = n3449 ^ n3309;
  assign n3444 = n3392 ^ n3385;
  assign n3445 = n3399 ^ n3385;
  assign n3446 = n3444 & ~n3445;
  assign n3447 = n3446 ^ n3392;
  assign n3451 = n3450 ^ n3447;
  assign n3456 = n3455 ^ n3451;
  assign n3440 = n3255 ^ n3247;
  assign n3441 = n3248 & n3440;
  assign n3442 = n3441 ^ n3245;
  assign n3432 = ~x5 & n2742;
  assign n3433 = ~x4 & n2746;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435 = x5 & n2749;
  assign n3436 = x4 & n2751;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = n3434 & n3437;
  assign n3439 = n3438 ^ x33;
  assign n3443 = n3442 ^ n3439;
  assign n3457 = n3456 ^ n3443;
  assign n3461 = n3460 ^ n3457;
  assign n3478 = n3477 ^ n3461;
  assign n3609 = n3608 ^ n3478;
  assign n3613 = n3612 ^ n3609;
  assign n3617 = n3616 ^ n3613;
  assign n3621 = n3620 ^ n3617;
  assign n3804 = n3620 ^ n3613;
  assign n3805 = n3617 & n3804;
  assign n3806 = n3805 ^ n3620;
  assign n3800 = n3612 ^ n3608;
  assign n3801 = ~n3609 & n3800;
  assign n3802 = n3801 ^ n3478;
  assign n3796 = n3607 ^ n3603;
  assign n3797 = n3604 & n3796;
  assign n3798 = n3797 ^ n3600;
  assign n3791 = n3472 ^ n3461;
  assign n3792 = ~n3477 & n3791;
  assign n3793 = n3792 ^ n3461;
  assign n3787 = n3599 ^ n3595;
  assign n3788 = ~n3596 & ~n3787;
  assign n3789 = n3788 ^ n3549;
  assign n3782 = n3460 ^ n3443;
  assign n3783 = n3460 ^ n3456;
  assign n3784 = n3782 & ~n3783;
  assign n3785 = n3784 ^ n3443;
  assign n3775 = n3563 ^ n3556;
  assign n3776 = n3570 ^ n3556;
  assign n3777 = n3775 & ~n3776;
  assign n3778 = n3777 ^ n3563;
  assign n3766 = x20 & n813;
  assign n3767 = x19 & n817;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = ~x20 & n820;
  assign n3770 = ~x19 & n822;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = n3768 & n3771;
  assign n3759 = ~x6 & n2742;
  assign n3760 = ~x5 & n2746;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = x6 & n2749;
  assign n3763 = x5 & n2751;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = n3761 & n3764;
  assign n3773 = n3772 ^ n3765;
  assign n3752 = ~x4 & n3163;
  assign n3753 = ~x3 & n3167;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = x4 & n3170;
  assign n3756 = x3 & n3172;
  assign n3757 = ~n3755 & ~n3756;
  assign n3758 = n3754 & n3757;
  assign n3774 = n3773 ^ n3758;
  assign n3779 = n3778 ^ n3774;
  assign n3743 = x16 & n1275;
  assign n3744 = x15 & n1279;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = ~x16 & n1282;
  assign n3747 = ~x15 & n1284;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = n3745 & n3748;
  assign n3736 = ~x18 & n1037;
  assign n3737 = ~x17 & n1041;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = x18 & n1044;
  assign n3740 = x17 & n1046;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = n3738 & n3741;
  assign n3750 = n3749 ^ n3742;
  assign n3729 = ~x24 & n460;
  assign n3730 = ~x23 & n462;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = x24 & n453;
  assign n3733 = x23 & n457;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = n3731 & n3734;
  assign n3751 = n3750 ^ n3735;
  assign n3780 = n3779 ^ n3751;
  assign n3718 = ~x14 & n1439;
  assign n3719 = ~x13 & n1443;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = x14 & n1446;
  assign n3722 = x13 & n1448;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = n3720 & n3723;
  assign n3711 = ~x12 & n1734;
  assign n3712 = ~x11 & n1738;
  assign n3713 = ~n3711 & ~n3712;
  assign n3714 = x12 & n1741;
  assign n3715 = x11 & n1743;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = n3713 & n3716;
  assign n3725 = n3724 ^ n3717;
  assign n3704 = ~x28 & n225;
  assign n3705 = ~x27 & n229;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = x28 & n232;
  assign n3708 = x27 & n234;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n3706 & n3709;
  assign n3726 = n3725 ^ n3710;
  assign n3695 = ~x30 & n159;
  assign n3696 = ~x29 & n163;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = x30 & n166;
  assign n3699 = x29 & n168;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = n3697 & n3700;
  assign n3688 = ~x26 & n344;
  assign n3689 = ~x25 & n348;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = x26 & n351;
  assign n3692 = x25 & n353;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = n3690 & n3693;
  assign n3702 = n3701 ^ n3694;
  assign n3687 = x2 & x63;
  assign n3703 = n3702 ^ n3687;
  assign n3727 = n3726 ^ n3703;
  assign n3678 = ~x10 & n2013;
  assign n3679 = ~x9 & n2017;
  assign n3680 = ~n3678 & ~n3679;
  assign n3681 = x10 & n2020;
  assign n3682 = x9 & n2022;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n3680 & n3683;
  assign n3671 = ~x22 & n618;
  assign n3672 = ~x21 & n622;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = x22 & n625;
  assign n3675 = x21 & n627;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = n3673 & n3676;
  assign n3685 = n3684 ^ n3677;
  assign n3664 = ~x8 & n2463;
  assign n3665 = ~x7 & n2465;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = x8 & n2456;
  assign n3668 = x7 & n2460;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = n3666 & n3669;
  assign n3686 = n3685 ^ n3670;
  assign n3728 = n3727 ^ n3686;
  assign n3781 = n3780 ^ n3728;
  assign n3786 = n3785 ^ n3781;
  assign n3790 = n3789 ^ n3786;
  assign n3794 = n3793 ^ n3790;
  assign n3658 = n3471 ^ n3464;
  assign n3659 = n3471 ^ n3467;
  assign n3660 = n3658 & ~n3659;
  assign n3661 = n3660 ^ n3464;
  assign n3653 = n3455 ^ n3447;
  assign n3654 = ~n3451 & n3653;
  assign n3655 = n3654 ^ n3455;
  assign n3650 = n3442 ^ n3438;
  assign n3651 = ~n3439 & n3650;
  assign n3652 = n3651 ^ x33;
  assign n3656 = n3655 ^ n3652;
  assign n3646 = n3515 ^ n3508;
  assign n3647 = ~n3523 & n3646;
  assign n3648 = n3647 ^ n3508;
  assign n3642 = n3538 ^ n3531;
  assign n3643 = ~n3546 & n3642;
  assign n3644 = n3643 ^ n3531;
  assign n3639 = n3499 ^ n3485;
  assign n3640 = n3500 & ~n3639;
  assign n3641 = n3640 ^ n3492;
  assign n3645 = n3644 ^ n3641;
  assign n3649 = n3648 ^ n3645;
  assign n3657 = n3656 ^ n3649;
  assign n3662 = n3661 ^ n3657;
  assign n3634 = n3524 ^ n3501;
  assign n3635 = n3547 ^ n3501;
  assign n3636 = n3634 & ~n3635;
  assign n3637 = n3636 ^ n3524;
  assign n3630 = n3589 ^ n3572;
  assign n3631 = n3594 & ~n3630;
  assign n3632 = n3631 ^ n3572;
  assign n3626 = n3580 ^ n3573;
  assign n3627 = ~n3588 & ~n3626;
  assign n3628 = n3627 ^ n3573;
  assign n3622 = x35 ^ x31;
  assign n3623 = n92 & n3622;
  assign n3624 = ~n89 & ~n3623;
  assign n3625 = n3624 ^ x33;
  assign n3629 = n3628 ^ n3625;
  assign n3633 = n3632 ^ n3629;
  assign n3638 = n3637 ^ n3633;
  assign n3663 = n3662 ^ n3638;
  assign n3795 = n3794 ^ n3663;
  assign n3799 = n3798 ^ n3795;
  assign n3803 = n3802 ^ n3799;
  assign n3807 = n3806 ^ n3803;
  assign n3988 = n3806 ^ n3799;
  assign n3989 = ~n3803 & ~n3988;
  assign n3990 = n3989 ^ n3806;
  assign n3984 = n3798 ^ n3794;
  assign n3985 = n3795 & n3984;
  assign n3986 = n3985 ^ n3663;
  assign n3979 = n3793 ^ n3786;
  assign n3980 = n3793 ^ n3789;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n3981 ^ n3786;
  assign n3974 = n3657 ^ n3638;
  assign n3975 = n3662 & ~n3974;
  assign n3976 = n3975 ^ n3638;
  assign n3970 = n3785 ^ n3780;
  assign n3971 = ~n3781 & ~n3970;
  assign n3972 = n3971 ^ n3728;
  assign n3965 = n3628 ^ n3624;
  assign n3966 = ~n3625 & ~n3965;
  assign n3967 = n3966 ^ x33;
  assign n3961 = n3648 ^ n3644;
  assign n3962 = n3645 & ~n3961;
  assign n3963 = n3962 ^ n3641;
  assign n3957 = n3694 ^ n3687;
  assign n3958 = ~n3702 & ~n3957;
  assign n3959 = n3958 ^ n3687;
  assign n3949 = x5 & n3170;
  assign n3950 = x4 & n3172;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = ~x5 & n3163;
  assign n3953 = ~x4 & n3167;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = n3951 & n3954;
  assign n3956 = n3955 ^ n3624;
  assign n3960 = n3959 ^ n3956;
  assign n3964 = n3963 ^ n3960;
  assign n3968 = n3967 ^ n3964;
  assign n3943 = n3765 ^ n3758;
  assign n3944 = ~n3773 & n3943;
  assign n3945 = n3944 ^ n3758;
  assign n3934 = ~x19 & n1037;
  assign n3935 = ~x18 & n1041;
  assign n3936 = ~n3934 & ~n3935;
  assign n3937 = x19 & n1044;
  assign n3938 = x18 & n1046;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = n3936 & n3939;
  assign n3933 = x3 & x63;
  assign n3941 = n3940 ^ n3933;
  assign n3926 = ~x17 & n1282;
  assign n3927 = ~x16 & n1284;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = x17 & n1275;
  assign n3930 = x16 & n1279;
  assign n3931 = ~n3929 & ~n3930;
  assign n3932 = n3928 & n3931;
  assign n3942 = n3941 ^ n3932;
  assign n3946 = n3945 ^ n3942;
  assign n3917 = x31 & n166;
  assign n3918 = x30 & n168;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~x31 & n159;
  assign n3921 = ~x30 & n163;
  assign n3922 = ~n3920 & ~n3921;
  assign n3923 = n3919 & n3922;
  assign n3916 = ~n89 & ~n93;
  assign n3924 = n3923 ^ n3916;
  assign n3909 = x27 & n351;
  assign n3910 = x26 & n353;
  assign n3911 = ~n3909 & ~n3910;
  assign n3912 = ~x27 & n344;
  assign n3913 = ~x26 & n348;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = n3911 & n3914;
  assign n3925 = n3924 ^ n3915;
  assign n3947 = n3946 ^ n3925;
  assign n3898 = ~x15 & n1439;
  assign n3899 = ~x14 & n1443;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = x15 & n1446;
  assign n3902 = x14 & n1448;
  assign n3903 = ~n3901 & ~n3902;
  assign n3904 = n3900 & n3903;
  assign n3891 = ~x25 & n460;
  assign n3892 = ~x24 & n462;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = x25 & n453;
  assign n3895 = x24 & n457;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = n3893 & n3896;
  assign n3905 = n3904 ^ n3897;
  assign n3884 = ~x13 & n1734;
  assign n3885 = ~x12 & n1738;
  assign n3886 = ~n3884 & ~n3885;
  assign n3887 = x13 & n1741;
  assign n3888 = x12 & n1743;
  assign n3889 = ~n3887 & ~n3888;
  assign n3890 = n3886 & n3889;
  assign n3906 = n3905 ^ n3890;
  assign n3875 = x9 & n2456;
  assign n3876 = x8 & n2460;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = ~x9 & n2463;
  assign n3879 = ~x8 & n2465;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = n3877 & n3880;
  assign n3868 = ~x21 & n820;
  assign n3869 = ~x20 & n822;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = x21 & n813;
  assign n3872 = x20 & n817;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = n3870 & n3873;
  assign n3882 = n3881 ^ n3874;
  assign n3861 = ~x7 & n2742;
  assign n3862 = ~x6 & n2746;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = x7 & n2749;
  assign n3865 = x6 & n2751;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = n3863 & n3866;
  assign n3883 = n3882 ^ n3867;
  assign n3907 = n3906 ^ n3883;
  assign n3852 = x23 & n625;
  assign n3853 = x22 & n627;
  assign n3854 = ~n3852 & ~n3853;
  assign n3855 = ~x23 & n618;
  assign n3856 = ~x22 & n622;
  assign n3857 = ~n3855 & ~n3856;
  assign n3858 = n3854 & n3857;
  assign n3845 = ~x29 & n225;
  assign n3846 = ~x28 & n229;
  assign n3847 = ~n3845 & ~n3846;
  assign n3848 = x29 & n232;
  assign n3849 = x28 & n234;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = n3847 & n3850;
  assign n3859 = n3858 ^ n3851;
  assign n3838 = x11 & n2020;
  assign n3839 = x10 & n2022;
  assign n3840 = ~n3838 & ~n3839;
  assign n3841 = ~x11 & n2013;
  assign n3842 = ~x10 & n2017;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = n3840 & n3843;
  assign n3860 = n3859 ^ n3844;
  assign n3908 = n3907 ^ n3860;
  assign n3948 = n3947 ^ n3908;
  assign n3969 = n3968 ^ n3948;
  assign n3973 = n3972 ^ n3969;
  assign n3977 = n3976 ^ n3973;
  assign n3833 = n3652 ^ n3649;
  assign n3834 = n3656 & ~n3833;
  assign n3835 = n3834 ^ n3649;
  assign n3829 = n3637 ^ n3629;
  assign n3830 = n3637 ^ n3632;
  assign n3831 = n3829 & ~n3830;
  assign n3832 = n3831 ^ n3629;
  assign n3836 = n3835 ^ n3832;
  assign n3824 = n3774 ^ n3751;
  assign n3825 = n3778 ^ n3751;
  assign n3826 = n3824 & ~n3825;
  assign n3827 = n3826 ^ n3774;
  assign n3819 = n3703 ^ n3686;
  assign n3820 = n3726 ^ n3686;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = n3821 ^ n3703;
  assign n3815 = n3684 ^ n3670;
  assign n3816 = n3685 & ~n3815;
  assign n3817 = n3816 ^ n3677;
  assign n3811 = n3749 ^ n3735;
  assign n3812 = n3750 & ~n3811;
  assign n3813 = n3812 ^ n3742;
  assign n3808 = n3717 ^ n3710;
  assign n3809 = ~n3725 & n3808;
  assign n3810 = n3809 ^ n3710;
  assign n3814 = n3813 ^ n3810;
  assign n3818 = n3817 ^ n3814;
  assign n3823 = n3822 ^ n3818;
  assign n3828 = n3827 ^ n3823;
  assign n3837 = n3836 ^ n3828;
  assign n3978 = n3977 ^ n3837;
  assign n3983 = n3982 ^ n3978;
  assign n3987 = n3986 ^ n3983;
  assign n3991 = n3990 ^ n3987;
  assign n4168 = n3990 ^ n3983;
  assign n4169 = n3987 & ~n4168;
  assign n4170 = n4169 ^ n3990;
  assign n4164 = n3982 ^ n3977;
  assign n4165 = ~n3978 & n4164;
  assign n4166 = n4165 ^ n3837;
  assign n4160 = n3976 ^ n3972;
  assign n4161 = n3973 & n4160;
  assign n4162 = n4161 ^ n3969;
  assign n4155 = n3832 ^ n3828;
  assign n4156 = ~n3836 & ~n4155;
  assign n4157 = n4156 ^ n3828;
  assign n4151 = n3968 ^ n3947;
  assign n4152 = n3948 & n4151;
  assign n4153 = n4152 ^ n3908;
  assign n4146 = n3967 ^ n3960;
  assign n4147 = n3967 ^ n3963;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = n4148 ^ n3960;
  assign n4142 = n3883 ^ n3860;
  assign n4143 = ~n3907 & n4142;
  assign n4144 = n4143 ^ n3860;
  assign n4131 = ~x24 & n618;
  assign n4132 = ~x23 & n622;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = x24 & n625;
  assign n4135 = x23 & n627;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = n4133 & n4136;
  assign n4124 = ~x16 & n1439;
  assign n4125 = ~x15 & n1443;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = x16 & n1446;
  assign n4128 = x15 & n1448;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = n4126 & n4129;
  assign n4138 = n4137 ^ n4130;
  assign n4117 = x14 & n1741;
  assign n4118 = x13 & n1743;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = ~x14 & n1734;
  assign n4121 = ~x13 & n1738;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = n4119 & n4122;
  assign n4139 = n4138 ^ n4123;
  assign n4108 = x8 & n2749;
  assign n4109 = x7 & n2751;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = ~x8 & n2742;
  assign n4112 = ~x7 & n2746;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = n4110 & n4113;
  assign n4101 = x10 & n2456;
  assign n4102 = x9 & n2460;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~x10 & n2463;
  assign n4105 = ~x9 & n2465;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = n4103 & n4106;
  assign n4115 = n4114 ^ n4107;
  assign n4094 = ~x20 & n1037;
  assign n4095 = ~x19 & n1041;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = x20 & n1044;
  assign n4098 = x19 & n1046;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = n4096 & n4099;
  assign n4116 = n4115 ^ n4100;
  assign n4140 = n4139 ^ n4116;
  assign n4085 = ~x12 & n2013;
  assign n4086 = ~x11 & n2017;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = x12 & n2020;
  assign n4089 = x11 & n2022;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n4087 & n4090;
  assign n4078 = ~x28 & n344;
  assign n4079 = ~x27 & n348;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = x28 & n351;
  assign n4082 = x27 & n353;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = n4080 & n4083;
  assign n4092 = n4091 ^ n4084;
  assign n4071 = x22 & n813;
  assign n4072 = x21 & n817;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = ~x22 & n820;
  assign n4075 = ~x21 & n822;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = n4073 & n4076;
  assign n4093 = n4092 ^ n4077;
  assign n4141 = n4140 ^ n4093;
  assign n4145 = n4144 ^ n4141;
  assign n4150 = n4149 ^ n4145;
  assign n4154 = n4153 ^ n4150;
  assign n4158 = n4157 ^ n4154;
  assign n4066 = n3827 ^ n3822;
  assign n4067 = ~n3823 & n4066;
  assign n4068 = n4067 ^ n3818;
  assign n4062 = n3959 ^ n3955;
  assign n4063 = n3956 & n4062;
  assign n4064 = n4063 ^ n3624;
  assign n4057 = n3817 ^ n3810;
  assign n4058 = n3817 ^ n3813;
  assign n4059 = n4057 & ~n4058;
  assign n4060 = n4059 ^ n3810;
  assign n4048 = x6 & n3170;
  assign n4049 = x5 & n3172;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = ~x6 & n3163;
  assign n4052 = ~x5 & n3167;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = n4050 & n4053;
  assign n4047 = x4 & x63;
  assign n4055 = n4054 ^ n4047;
  assign n4044 = x37 ^ x31;
  assign n4045 = n162 & n4044;
  assign n4046 = ~n159 & ~n4045;
  assign n4056 = n4055 ^ n4046;
  assign n4061 = n4060 ^ n4056;
  assign n4065 = n4064 ^ n4061;
  assign n4069 = n4068 ^ n4065;
  assign n4038 = n3942 ^ n3925;
  assign n4039 = n3945 ^ n3925;
  assign n4040 = n4038 & n4039;
  assign n4041 = n4040 ^ n3942;
  assign n4033 = n3897 ^ n3890;
  assign n4034 = n3904 ^ n3890;
  assign n4035 = n4033 & ~n4034;
  assign n4036 = n4035 ^ n3897;
  assign n4028 = n3933 ^ n3932;
  assign n4029 = n3940 ^ n3932;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n4030 ^ n3933;
  assign n4024 = n3916 ^ n3915;
  assign n4025 = n3923 ^ n3915;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = n4026 ^ n3916;
  assign n4032 = n4031 ^ n4027;
  assign n4037 = n4036 ^ n4032;
  assign n4042 = n4041 ^ n4037;
  assign n4018 = n3874 ^ n3867;
  assign n4019 = n3881 ^ n3867;
  assign n4020 = n4018 & ~n4019;
  assign n4021 = n4020 ^ n3874;
  assign n4015 = n3858 ^ n3844;
  assign n4016 = n3859 & ~n4015;
  assign n4017 = n4016 ^ n3851;
  assign n4022 = n4021 ^ n4017;
  assign n4006 = ~x30 & n225;
  assign n4007 = ~x29 & n229;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = x30 & n232;
  assign n4010 = x29 & n234;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = n4008 & n4011;
  assign n3999 = ~x26 & n460;
  assign n4000 = ~x25 & n462;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = x26 & n453;
  assign n4003 = x25 & n457;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = n4001 & n4004;
  assign n4013 = n4012 ^ n4005;
  assign n3992 = x18 & n1275;
  assign n3993 = x17 & n1279;
  assign n3994 = ~n3992 & ~n3993;
  assign n3995 = ~x18 & n1282;
  assign n3996 = ~x17 & n1284;
  assign n3997 = ~n3995 & ~n3996;
  assign n3998 = n3994 & n3997;
  assign n4014 = n4013 ^ n3998;
  assign n4023 = n4022 ^ n4014;
  assign n4043 = n4042 ^ n4023;
  assign n4070 = n4069 ^ n4043;
  assign n4159 = n4158 ^ n4070;
  assign n4163 = n4162 ^ n4159;
  assign n4167 = n4166 ^ n4163;
  assign n4171 = n4170 ^ n4167;
  assign n4342 = n4170 ^ n4163;
  assign n4343 = n4167 & ~n4342;
  assign n4344 = n4343 ^ n4170;
  assign n4338 = n4162 ^ n4158;
  assign n4339 = ~n4159 & n4338;
  assign n4340 = n4339 ^ n4070;
  assign n4334 = n4157 ^ n4153;
  assign n4335 = ~n4154 & n4334;
  assign n4336 = n4335 ^ n4150;
  assign n4328 = n4065 ^ n4043;
  assign n4329 = n4068 ^ n4043;
  assign n4330 = ~n4328 & n4329;
  assign n4331 = n4330 ^ n4065;
  assign n4324 = n4149 ^ n4144;
  assign n4325 = n4145 & n4324;
  assign n4326 = n4325 ^ n4141;
  assign n4318 = n4036 ^ n4027;
  assign n4319 = n4036 ^ n4031;
  assign n4320 = ~n4318 & n4319;
  assign n4321 = n4320 ^ n4027;
  assign n4313 = n4047 ^ n4046;
  assign n4314 = n4054 ^ n4046;
  assign n4315 = n4313 & n4314;
  assign n4316 = n4315 ^ n4047;
  assign n4304 = x13 & n2020;
  assign n4305 = x12 & n2022;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = ~x13 & n2013;
  assign n4308 = ~x12 & n2017;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = n4306 & n4309;
  assign n4297 = ~x15 & n1734;
  assign n4298 = ~x14 & n1738;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = x15 & n1741;
  assign n4301 = x14 & n1743;
  assign n4302 = ~n4300 & ~n4301;
  assign n4303 = n4299 & n4302;
  assign n4311 = n4310 ^ n4303;
  assign n4290 = ~x29 & n344;
  assign n4291 = ~x28 & n348;
  assign n4292 = ~n4290 & ~n4291;
  assign n4293 = x29 & n351;
  assign n4294 = x28 & n353;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = n4292 & n4295;
  assign n4312 = n4311 ^ n4296;
  assign n4317 = n4316 ^ n4312;
  assign n4322 = n4321 ^ n4317;
  assign n4285 = n4116 ^ n4093;
  assign n4286 = n4139 ^ n4093;
  assign n4287 = n4285 & ~n4286;
  assign n4288 = n4287 ^ n4116;
  assign n4274 = ~x7 & n3163;
  assign n4275 = ~x6 & n3167;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = x7 & n3170;
  assign n4278 = x6 & n3172;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = n4276 & n4279;
  assign n4267 = ~x21 & n1037;
  assign n4268 = ~x20 & n1041;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = x21 & n1044;
  assign n4271 = x20 & n1046;
  assign n4272 = ~n4270 & ~n4271;
  assign n4273 = n4269 & n4272;
  assign n4281 = n4280 ^ n4273;
  assign n4266 = x5 & x63;
  assign n4282 = n4281 ^ n4266;
  assign n4257 = ~x31 & n225;
  assign n4258 = ~x30 & n229;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = x31 & n232;
  assign n4261 = x30 & n234;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = n4259 & n4262;
  assign n4256 = ~n159 & ~n163;
  assign n4264 = n4263 ^ n4256;
  assign n4249 = ~x27 & n460;
  assign n4250 = ~x26 & n462;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = x27 & n453;
  assign n4253 = x26 & n457;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = n4251 & n4254;
  assign n4265 = n4264 ^ n4255;
  assign n4283 = n4282 ^ n4265;
  assign n4240 = ~x11 & n2463;
  assign n4241 = ~x10 & n2465;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = x11 & n2456;
  assign n4244 = x10 & n2460;
  assign n4245 = ~n4243 & ~n4244;
  assign n4246 = n4242 & n4245;
  assign n4233 = ~x23 & n820;
  assign n4234 = ~x22 & n822;
  assign n4235 = ~n4233 & ~n4234;
  assign n4236 = x23 & n813;
  assign n4237 = x22 & n817;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = n4235 & n4238;
  assign n4247 = n4246 ^ n4239;
  assign n4226 = ~x9 & n2742;
  assign n4227 = ~x8 & n2746;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = x9 & n2749;
  assign n4230 = x8 & n2751;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = n4228 & n4231;
  assign n4248 = n4247 ^ n4232;
  assign n4284 = n4283 ^ n4248;
  assign n4289 = n4288 ^ n4284;
  assign n4323 = n4322 ^ n4289;
  assign n4327 = n4326 ^ n4323;
  assign n4332 = n4331 ^ n4327;
  assign n4221 = n4037 ^ n4023;
  assign n4222 = n4042 & n4221;
  assign n4223 = n4222 ^ n4023;
  assign n4217 = n4064 ^ n4056;
  assign n4218 = n4064 ^ n4060;
  assign n4219 = n4217 & ~n4218;
  assign n4220 = n4219 ^ n4056;
  assign n4224 = n4223 ^ n4220;
  assign n4213 = n4017 ^ n4014;
  assign n4214 = ~n4022 & n4213;
  assign n4215 = n4214 ^ n4014;
  assign n4208 = n4137 ^ n4123;
  assign n4209 = n4138 & ~n4208;
  assign n4210 = n4209 ^ n4130;
  assign n4204 = n4012 ^ n3998;
  assign n4205 = n4013 & ~n4204;
  assign n4206 = n4205 ^ n4005;
  assign n4207 = n4206 ^ n4046;
  assign n4211 = n4210 ^ n4207;
  assign n4198 = n4084 ^ n4077;
  assign n4199 = n4091 ^ n4077;
  assign n4200 = n4198 & ~n4199;
  assign n4201 = n4200 ^ n4084;
  assign n4195 = n4107 ^ n4100;
  assign n4196 = ~n4115 & n4195;
  assign n4197 = n4196 ^ n4100;
  assign n4202 = n4201 ^ n4197;
  assign n4186 = x17 & n1446;
  assign n4187 = x16 & n1448;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~x17 & n1439;
  assign n4190 = ~x16 & n1443;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = n4188 & n4191;
  assign n4179 = ~x19 & n1282;
  assign n4180 = ~x18 & n1284;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = x19 & n1275;
  assign n4183 = x18 & n1279;
  assign n4184 = ~n4182 & ~n4183;
  assign n4185 = n4181 & n4184;
  assign n4193 = n4192 ^ n4185;
  assign n4172 = ~x25 & n618;
  assign n4173 = ~x24 & n622;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = x25 & n625;
  assign n4176 = x24 & n627;
  assign n4177 = ~n4175 & ~n4176;
  assign n4178 = n4174 & n4177;
  assign n4194 = n4193 ^ n4178;
  assign n4203 = n4202 ^ n4194;
  assign n4212 = n4211 ^ n4203;
  assign n4216 = n4215 ^ n4212;
  assign n4225 = n4224 ^ n4216;
  assign n4333 = n4332 ^ n4225;
  assign n4337 = n4336 ^ n4333;
  assign n4341 = n4340 ^ n4337;
  assign n4345 = n4344 ^ n4341;
  assign n4505 = n4344 ^ n4337;
  assign n4506 = ~n4341 & n4505;
  assign n4507 = n4506 ^ n4344;
  assign n4501 = n4336 ^ n4332;
  assign n4502 = n4333 & n4501;
  assign n4503 = n4502 ^ n4225;
  assign n4497 = n4331 ^ n4326;
  assign n4498 = n4327 & ~n4497;
  assign n4499 = n4498 ^ n4323;
  assign n4493 = n4220 ^ n4216;
  assign n4494 = ~n4224 & n4493;
  assign n4495 = n4494 ^ n4216;
  assign n4488 = n4322 ^ n4288;
  assign n4489 = n4289 & ~n4488;
  assign n4490 = n4489 ^ n4284;
  assign n4484 = n4321 ^ n4316;
  assign n4485 = ~n4317 & ~n4484;
  assign n4486 = n4485 ^ n4312;
  assign n4479 = n4265 ^ n4248;
  assign n4480 = n4282 ^ n4248;
  assign n4481 = ~n4479 & n4480;
  assign n4482 = n4481 ^ n4265;
  assign n4474 = n4273 ^ n4266;
  assign n4475 = ~n4281 & ~n4474;
  assign n4476 = n4475 ^ n4266;
  assign n4465 = ~x8 & n3163;
  assign n4466 = ~x7 & n3167;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = x8 & n3170;
  assign n4469 = x7 & n3172;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = n4467 & n4470;
  assign n4458 = ~x28 & n460;
  assign n4459 = ~x27 & n462;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = x28 & n453;
  assign n4462 = x27 & n457;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = n4460 & n4463;
  assign n4472 = n4471 ^ n4464;
  assign n4457 = x6 & x63;
  assign n4473 = n4472 ^ n4457;
  assign n4477 = n4476 ^ n4473;
  assign n4448 = ~x18 & n1439;
  assign n4449 = ~x17 & n1443;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = x18 & n1446;
  assign n4452 = x17 & n1448;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = n4450 & n4453;
  assign n4441 = ~x26 & n618;
  assign n4442 = ~x25 & n622;
  assign n4443 = ~n4441 & ~n4442;
  assign n4444 = x26 & n625;
  assign n4445 = x25 & n627;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = n4443 & n4446;
  assign n4455 = n4454 ^ n4447;
  assign n4434 = ~x16 & n1734;
  assign n4435 = ~x15 & n1738;
  assign n4436 = ~n4434 & ~n4435;
  assign n4437 = x16 & n1741;
  assign n4438 = x15 & n1743;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = n4436 & n4439;
  assign n4456 = n4455 ^ n4440;
  assign n4478 = n4477 ^ n4456;
  assign n4483 = n4482 ^ n4478;
  assign n4487 = n4486 ^ n4483;
  assign n4491 = n4490 ^ n4487;
  assign n4429 = n4215 ^ n4211;
  assign n4430 = n4212 & ~n4429;
  assign n4431 = n4430 ^ n4203;
  assign n4424 = n4239 ^ n4232;
  assign n4425 = ~n4247 & n4424;
  assign n4426 = n4425 ^ n4232;
  assign n4416 = ~x20 & n1282;
  assign n4417 = ~x19 & n1284;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = x20 & n1275;
  assign n4420 = x19 & n1279;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = n4418 & n4421;
  assign n4409 = ~x30 & n344;
  assign n4410 = ~x29 & n348;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = x30 & n351;
  assign n4413 = x29 & n353;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = n4411 & n4414;
  assign n4423 = n4422 ^ n4415;
  assign n4427 = n4426 ^ n4423;
  assign n4399 = ~x14 & n2013;
  assign n4400 = ~x13 & n2017;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = x14 & n2020;
  assign n4403 = x13 & n2022;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = n4401 & n4404;
  assign n4392 = ~x24 & n820;
  assign n4393 = ~x23 & n822;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = x24 & n813;
  assign n4396 = x23 & n817;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = n4394 & n4397;
  assign n4406 = n4405 ^ n4398;
  assign n4385 = x12 & n2456;
  assign n4386 = x11 & n2460;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = ~x12 & n2463;
  assign n4389 = ~x11 & n2465;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = n4387 & n4390;
  assign n4407 = n4406 ^ n4391;
  assign n4376 = ~x22 & n1037;
  assign n4377 = ~x21 & n1041;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = x22 & n1044;
  assign n4380 = x21 & n1046;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = n4378 & n4381;
  assign n4373 = x39 ^ x31;
  assign n4374 = n228 & n4373;
  assign n4375 = ~n225 & ~n4374;
  assign n4383 = n4382 ^ n4375;
  assign n4366 = ~x10 & n2742;
  assign n4367 = ~x9 & n2746;
  assign n4368 = ~n4366 & ~n4367;
  assign n4369 = x10 & n2749;
  assign n4370 = x9 & n2751;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = n4368 & n4371;
  assign n4384 = n4383 ^ n4372;
  assign n4408 = n4407 ^ n4384;
  assign n4428 = n4427 ^ n4408;
  assign n4432 = n4431 ^ n4428;
  assign n4362 = n4197 ^ n4194;
  assign n4363 = ~n4202 & n4362;
  assign n4364 = n4363 ^ n4194;
  assign n4358 = n4210 ^ n4206;
  assign n4359 = n4207 & ~n4358;
  assign n4360 = n4359 ^ n4046;
  assign n4354 = n4310 ^ n4296;
  assign n4355 = n4311 & ~n4354;
  assign n4356 = n4355 ^ n4303;
  assign n4350 = n4185 ^ n4178;
  assign n4351 = ~n4193 & n4350;
  assign n4352 = n4351 ^ n4178;
  assign n4346 = n4256 ^ n4255;
  assign n4347 = n4263 ^ n4255;
  assign n4348 = ~n4346 & ~n4347;
  assign n4349 = n4348 ^ n4256;
  assign n4353 = n4352 ^ n4349;
  assign n4357 = n4356 ^ n4353;
  assign n4361 = n4360 ^ n4357;
  assign n4365 = n4364 ^ n4361;
  assign n4433 = n4432 ^ n4365;
  assign n4492 = n4491 ^ n4433;
  assign n4496 = n4495 ^ n4492;
  assign n4500 = n4499 ^ n4496;
  assign n4504 = n4503 ^ n4500;
  assign n4508 = n4507 ^ n4504;
  assign n4664 = n4507 ^ n4500;
  assign n4665 = n4504 & n4664;
  assign n4666 = n4665 ^ n4507;
  assign n4660 = n4499 ^ n4495;
  assign n4661 = ~n4496 & ~n4660;
  assign n4662 = n4661 ^ n4492;
  assign n4655 = n4487 ^ n4433;
  assign n4656 = n4490 ^ n4433;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = n4657 ^ n4487;
  assign n4650 = n4428 ^ n4365;
  assign n4651 = n4431 ^ n4365;
  assign n4652 = n4650 & n4651;
  assign n4653 = n4652 ^ n4428;
  assign n4645 = n4486 ^ n4482;
  assign n4646 = ~n4483 & n4645;
  assign n4647 = n4646 ^ n4478;
  assign n4640 = n4473 ^ n4456;
  assign n4641 = ~n4477 & ~n4640;
  assign n4642 = n4641 ^ n4456;
  assign n4635 = n4464 ^ n4457;
  assign n4636 = ~n4472 & ~n4635;
  assign n4637 = n4636 ^ n4457;
  assign n4626 = ~x17 & n1734;
  assign n4627 = ~x16 & n1738;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = x17 & n1741;
  assign n4630 = x16 & n1743;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = n4628 & n4631;
  assign n4619 = ~x19 & n1439;
  assign n4620 = ~x18 & n1443;
  assign n4621 = ~n4619 & ~n4620;
  assign n4622 = x19 & n1446;
  assign n4623 = x18 & n1448;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = n4621 & n4624;
  assign n4633 = n4632 ^ n4625;
  assign n4612 = ~x25 & n820;
  assign n4613 = ~x24 & n822;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = x25 & n813;
  assign n4616 = x24 & n817;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = n4614 & n4617;
  assign n4634 = n4633 ^ n4618;
  assign n4638 = n4637 ^ n4634;
  assign n4603 = ~x31 & n344;
  assign n4604 = ~x30 & n348;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = x31 & n351;
  assign n4607 = x30 & n353;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = n4605 & n4608;
  assign n4602 = ~n225 & ~n229;
  assign n4610 = n4609 ^ n4602;
  assign n4595 = x27 & n625;
  assign n4596 = x26 & n627;
  assign n4597 = ~n4595 & ~n4596;
  assign n4598 = ~x27 & n618;
  assign n4599 = ~x26 & n622;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = n4597 & n4600;
  assign n4611 = n4610 ^ n4601;
  assign n4639 = n4638 ^ n4611;
  assign n4643 = n4642 ^ n4639;
  assign n4584 = ~x13 & n2463;
  assign n4585 = ~x12 & n2465;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = x13 & n2456;
  assign n4588 = x12 & n2460;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = n4586 & n4589;
  assign n4577 = x15 & n2020;
  assign n4578 = x14 & n2022;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = ~x15 & n2013;
  assign n4581 = ~x14 & n2017;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = n4579 & n4582;
  assign n4591 = n4590 ^ n4583;
  assign n4570 = ~x29 & n460;
  assign n4571 = ~x28 & n462;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = x29 & n453;
  assign n4574 = x28 & n457;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = n4572 & n4575;
  assign n4592 = n4591 ^ n4576;
  assign n4561 = ~x11 & n2742;
  assign n4562 = ~x10 & n2746;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = x11 & n2749;
  assign n4565 = x10 & n2751;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4563 & n4566;
  assign n4554 = x23 & n1044;
  assign n4555 = x22 & n1046;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = ~x23 & n1037;
  assign n4558 = ~x22 & n1041;
  assign n4559 = ~n4557 & ~n4558;
  assign n4560 = n4556 & n4559;
  assign n4568 = n4567 ^ n4560;
  assign n4547 = x9 & n3170;
  assign n4548 = x8 & n3172;
  assign n4549 = ~n4547 & ~n4548;
  assign n4550 = ~x9 & n3163;
  assign n4551 = ~x8 & n3167;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = n4549 & n4552;
  assign n4569 = n4568 ^ n4553;
  assign n4593 = n4592 ^ n4569;
  assign n4538 = ~x21 & n1282;
  assign n4539 = ~x20 & n1284;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = x21 & n1275;
  assign n4542 = x20 & n1279;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = n4540 & n4543;
  assign n4537 = x7 & x63;
  assign n4545 = n4544 ^ n4537;
  assign n4546 = n4545 ^ n4415;
  assign n4594 = n4593 ^ n4546;
  assign n4644 = n4643 ^ n4594;
  assign n4648 = n4647 ^ n4644;
  assign n4532 = n4364 ^ n4357;
  assign n4533 = n4364 ^ n4360;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = n4534 ^ n4357;
  assign n4528 = n4427 ^ n4407;
  assign n4529 = n4408 & n4528;
  assign n4530 = n4529 ^ n4384;
  assign n4523 = n4356 ^ n4352;
  assign n4524 = ~n4353 & ~n4523;
  assign n4525 = n4524 ^ n4349;
  assign n4520 = n4426 ^ n4422;
  assign n4521 = ~n4423 & ~n4520;
  assign n4522 = n4521 ^ n4415;
  assign n4526 = n4525 ^ n4522;
  assign n4516 = n4382 ^ n4372;
  assign n4517 = n4383 & ~n4516;
  assign n4518 = n4517 ^ n4375;
  assign n4512 = n4447 ^ n4440;
  assign n4513 = ~n4455 & n4512;
  assign n4514 = n4513 ^ n4440;
  assign n4509 = n4398 ^ n4391;
  assign n4510 = ~n4406 & n4509;
  assign n4511 = n4510 ^ n4391;
  assign n4515 = n4514 ^ n4511;
  assign n4519 = n4518 ^ n4515;
  assign n4527 = n4526 ^ n4519;
  assign n4531 = n4530 ^ n4527;
  assign n4536 = n4535 ^ n4531;
  assign n4649 = n4648 ^ n4536;
  assign n4654 = n4653 ^ n4649;
  assign n4659 = n4658 ^ n4654;
  assign n4663 = n4662 ^ n4659;
  assign n4667 = n4666 ^ n4663;
  assign n4816 = n4666 ^ n4659;
  assign n4817 = n4663 & ~n4816;
  assign n4818 = n4817 ^ n4666;
  assign n4811 = n4658 ^ n4653;
  assign n4812 = n4658 ^ n4649;
  assign n4813 = n4811 & n4812;
  assign n4814 = n4813 ^ n4653;
  assign n4806 = n4644 ^ n4536;
  assign n4807 = n4647 ^ n4536;
  assign n4808 = n4806 & n4807;
  assign n4809 = n4808 ^ n4644;
  assign n4801 = n4535 ^ n4527;
  assign n4802 = n4531 & n4801;
  assign n4803 = n4802 ^ n4530;
  assign n4797 = n4639 ^ n4594;
  assign n4798 = ~n4643 & ~n4797;
  assign n4799 = n4798 ^ n4594;
  assign n4793 = n4569 ^ n4546;
  assign n4794 = ~n4593 & ~n4793;
  assign n4795 = n4794 ^ n4546;
  assign n4789 = n4634 ^ n4611;
  assign n4790 = n4638 & ~n4789;
  assign n4791 = n4790 ^ n4611;
  assign n4784 = n4567 ^ n4553;
  assign n4785 = n4568 & ~n4784;
  assign n4786 = n4785 ^ n4560;
  assign n4780 = n4602 ^ n4601;
  assign n4781 = n4609 ^ n4601;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = n4782 ^ n4602;
  assign n4787 = n4786 ^ n4783;
  assign n4771 = x28 & n625;
  assign n4772 = x27 & n627;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~x28 & n618;
  assign n4775 = ~x27 & n622;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = n4773 & n4776;
  assign n4770 = x8 & x63;
  assign n4778 = n4777 ^ n4770;
  assign n4763 = ~x20 & n1439;
  assign n4764 = ~x19 & n1443;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = x20 & n1446;
  assign n4767 = x19 & n1448;
  assign n4768 = ~n4766 & ~n4767;
  assign n4769 = n4765 & n4768;
  assign n4779 = n4778 ^ n4769;
  assign n4788 = n4787 ^ n4779;
  assign n4792 = n4791 ^ n4788;
  assign n4796 = n4795 ^ n4792;
  assign n4800 = n4799 ^ n4796;
  assign n4804 = n4803 ^ n4800;
  assign n4758 = n4522 ^ n4519;
  assign n4759 = ~n4526 & ~n4758;
  assign n4760 = n4759 ^ n4519;
  assign n4747 = x22 & n1275;
  assign n4748 = x21 & n1279;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = ~x22 & n1282;
  assign n4751 = ~x21 & n1284;
  assign n4752 = ~n4750 & ~n4751;
  assign n4753 = n4749 & n4752;
  assign n4744 = x41 ^ x31;
  assign n4745 = n347 & n4744;
  assign n4746 = ~n344 & ~n4745;
  assign n4754 = n4753 ^ n4746;
  assign n4737 = ~x10 & n3163;
  assign n4738 = ~x9 & n3167;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = x10 & n3170;
  assign n4741 = x9 & n3172;
  assign n4742 = ~n4740 & ~n4741;
  assign n4743 = n4739 & n4742;
  assign n4755 = n4754 ^ n4743;
  assign n4728 = x26 & n813;
  assign n4729 = x25 & n817;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = ~x26 & n820;
  assign n4732 = ~x25 & n822;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = n4730 & n4733;
  assign n4721 = ~x18 & n1734;
  assign n4722 = ~x17 & n1738;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = x18 & n1741;
  assign n4725 = x17 & n1743;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = n4723 & n4726;
  assign n4735 = n4734 ^ n4727;
  assign n4714 = ~x16 & n2013;
  assign n4715 = ~x15 & n2017;
  assign n4716 = ~n4714 & ~n4715;
  assign n4717 = x16 & n2020;
  assign n4718 = x15 & n2022;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = n4716 & n4719;
  assign n4736 = n4735 ^ n4720;
  assign n4756 = n4755 ^ n4736;
  assign n4705 = ~x14 & n2463;
  assign n4706 = ~x13 & n2465;
  assign n4707 = ~n4705 & ~n4706;
  assign n4708 = x14 & n2456;
  assign n4709 = x13 & n2460;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = n4707 & n4710;
  assign n4698 = ~x24 & n1037;
  assign n4699 = ~x23 & n1041;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = x24 & n1044;
  assign n4702 = x23 & n1046;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = n4700 & n4703;
  assign n4712 = n4711 ^ n4704;
  assign n4691 = ~x12 & n2742;
  assign n4692 = ~x11 & n2746;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = x12 & n2749;
  assign n4695 = x11 & n2751;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = n4693 & n4696;
  assign n4713 = n4712 ^ n4697;
  assign n4757 = n4756 ^ n4713;
  assign n4761 = n4760 ^ n4757;
  assign n4686 = n4518 ^ n4514;
  assign n4687 = n4515 & ~n4686;
  assign n4688 = n4687 ^ n4511;
  assign n4683 = n4544 ^ n4415;
  assign n4684 = ~n4545 & ~n4683;
  assign n4685 = n4684 ^ n4537;
  assign n4689 = n4688 ^ n4685;
  assign n4679 = n4583 ^ n4576;
  assign n4680 = ~n4591 & n4679;
  assign n4681 = n4680 ^ n4576;
  assign n4675 = n4625 ^ n4618;
  assign n4676 = ~n4633 & n4675;
  assign n4677 = n4676 ^ n4618;
  assign n4668 = ~x30 & n460;
  assign n4669 = ~x29 & n462;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = x30 & n453;
  assign n4672 = x29 & n457;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n4670 & n4673;
  assign n4678 = n4677 ^ n4674;
  assign n4682 = n4681 ^ n4678;
  assign n4690 = n4689 ^ n4682;
  assign n4762 = n4761 ^ n4690;
  assign n4805 = n4804 ^ n4762;
  assign n4810 = n4809 ^ n4805;
  assign n4815 = n4814 ^ n4810;
  assign n4819 = n4818 ^ n4815;
  assign n4966 = n4818 ^ n4810;
  assign n4967 = n4815 & ~n4966;
  assign n4968 = n4967 ^ n4818;
  assign n4962 = n4809 ^ n4804;
  assign n4963 = ~n4805 & ~n4962;
  assign n4964 = n4963 ^ n4762;
  assign n4958 = n4803 ^ n4799;
  assign n4959 = ~n4800 & n4958;
  assign n4960 = n4959 ^ n4796;
  assign n4952 = n4757 ^ n4690;
  assign n4953 = n4760 ^ n4690;
  assign n4954 = n4952 & ~n4953;
  assign n4955 = n4954 ^ n4757;
  assign n4947 = n4795 ^ n4788;
  assign n4948 = n4795 ^ n4791;
  assign n4949 = ~n4947 & ~n4948;
  assign n4950 = n4949 ^ n4788;
  assign n4942 = n4736 ^ n4713;
  assign n4943 = n4755 ^ n4713;
  assign n4944 = n4942 & ~n4943;
  assign n4945 = n4944 ^ n4736;
  assign n4938 = n4783 ^ n4779;
  assign n4939 = n4787 & n4938;
  assign n4940 = n4939 ^ n4779;
  assign n4933 = n4727 ^ n4720;
  assign n4934 = n4734 ^ n4720;
  assign n4935 = n4933 & ~n4934;
  assign n4936 = n4935 ^ n4727;
  assign n4928 = n4746 ^ n4743;
  assign n4929 = n4753 ^ n4743;
  assign n4930 = n4928 & ~n4929;
  assign n4931 = n4930 ^ n4746;
  assign n4925 = n4777 ^ n4769;
  assign n4926 = ~n4778 & ~n4925;
  assign n4927 = n4926 ^ n4770;
  assign n4932 = n4931 ^ n4927;
  assign n4937 = n4936 ^ n4932;
  assign n4941 = n4940 ^ n4937;
  assign n4946 = n4945 ^ n4941;
  assign n4951 = n4950 ^ n4946;
  assign n4956 = n4955 ^ n4951;
  assign n4919 = n4685 ^ n4682;
  assign n4920 = n4688 ^ n4682;
  assign n4921 = n4919 & n4920;
  assign n4922 = n4921 ^ n4685;
  assign n4908 = ~x13 & n2742;
  assign n4909 = ~x12 & n2746;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = x13 & n2749;
  assign n4912 = x12 & n2751;
  assign n4913 = ~n4911 & ~n4912;
  assign n4914 = n4910 & n4913;
  assign n4901 = ~x15 & n2463;
  assign n4902 = ~x14 & n2465;
  assign n4903 = ~n4901 & ~n4902;
  assign n4904 = x15 & n2456;
  assign n4905 = x14 & n2460;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = n4903 & n4906;
  assign n4915 = n4914 ^ n4907;
  assign n4894 = ~x29 & n618;
  assign n4895 = ~x28 & n622;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = x29 & n625;
  assign n4898 = x28 & n627;
  assign n4899 = ~n4897 & ~n4898;
  assign n4900 = n4896 & n4899;
  assign n4916 = n4915 ^ n4900;
  assign n4885 = ~x31 & n460;
  assign n4886 = ~x30 & n462;
  assign n4887 = ~n4885 & ~n4886;
  assign n4888 = x31 & n453;
  assign n4889 = x30 & n457;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n4887 & n4890;
  assign n4884 = ~n344 & ~n348;
  assign n4892 = n4891 ^ n4884;
  assign n4877 = x27 & n813;
  assign n4878 = x26 & n817;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~x27 & n820;
  assign n4881 = ~x26 & n822;
  assign n4882 = ~n4880 & ~n4881;
  assign n4883 = n4879 & n4882;
  assign n4893 = n4892 ^ n4883;
  assign n4917 = n4916 ^ n4893;
  assign n4868 = ~x17 & n2013;
  assign n4869 = ~x16 & n2017;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = x17 & n2020;
  assign n4872 = x16 & n2022;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = n4870 & n4873;
  assign n4861 = x19 & n1741;
  assign n4862 = x18 & n1743;
  assign n4863 = ~n4861 & ~n4862;
  assign n4864 = ~x19 & n1734;
  assign n4865 = ~x18 & n1738;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = n4863 & n4866;
  assign n4875 = n4874 ^ n4867;
  assign n4854 = x25 & n1044;
  assign n4855 = x24 & n1046;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = ~x25 & n1037;
  assign n4858 = ~x24 & n1041;
  assign n4859 = ~n4857 & ~n4858;
  assign n4860 = n4856 & n4859;
  assign n4876 = n4875 ^ n4860;
  assign n4918 = n4917 ^ n4876;
  assign n4923 = n4922 ^ n4918;
  assign n4850 = n4681 ^ n4677;
  assign n4851 = ~n4678 & ~n4850;
  assign n4852 = n4851 ^ n4674;
  assign n4845 = n4704 ^ n4697;
  assign n4846 = ~n4712 & n4845;
  assign n4847 = n4846 ^ n4697;
  assign n4837 = ~x21 & n1439;
  assign n4838 = ~x20 & n1443;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = x21 & n1446;
  assign n4841 = x20 & n1448;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = n4839 & n4842;
  assign n4844 = n4843 ^ n4674;
  assign n4848 = n4847 ^ n4844;
  assign n4828 = ~x11 & n3163;
  assign n4829 = ~x10 & n3167;
  assign n4830 = ~n4828 & ~n4829;
  assign n4831 = x11 & n3170;
  assign n4832 = x10 & n3172;
  assign n4833 = ~n4831 & ~n4832;
  assign n4834 = n4830 & n4833;
  assign n4821 = ~x23 & n1282;
  assign n4822 = ~x22 & n1284;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = x23 & n1275;
  assign n4825 = x22 & n1279;
  assign n4826 = ~n4824 & ~n4825;
  assign n4827 = n4823 & n4826;
  assign n4835 = n4834 ^ n4827;
  assign n4820 = x9 & x63;
  assign n4836 = n4835 ^ n4820;
  assign n4849 = n4848 ^ n4836;
  assign n4853 = n4852 ^ n4849;
  assign n4924 = n4923 ^ n4853;
  assign n4957 = n4956 ^ n4924;
  assign n4961 = n4960 ^ n4957;
  assign n4965 = n4964 ^ n4961;
  assign n4969 = n4968 ^ n4965;
  assign n5105 = n4968 ^ n4961;
  assign n5106 = ~n4965 & ~n5105;
  assign n5107 = n5106 ^ n4968;
  assign n5101 = n4960 ^ n4956;
  assign n5102 = n4957 & ~n5101;
  assign n5103 = n5102 ^ n4924;
  assign n5097 = n4955 ^ n4950;
  assign n5098 = n4951 & ~n5097;
  assign n5099 = n5098 ^ n4946;
  assign n5091 = n4918 ^ n4853;
  assign n5092 = n4922 ^ n4853;
  assign n5093 = ~n5091 & n5092;
  assign n5094 = n5093 ^ n4918;
  assign n5087 = n4945 ^ n4937;
  assign n5088 = ~n4941 & ~n5087;
  assign n5089 = n5088 ^ n4945;
  assign n5083 = n4916 ^ n4876;
  assign n5084 = ~n4917 & ~n5083;
  assign n5085 = n5084 ^ n4893;
  assign n5079 = n4847 ^ n4843;
  assign n5080 = n4844 & ~n5079;
  assign n5081 = n5080 ^ n4674;
  assign n5075 = n4891 ^ n4883;
  assign n5076 = ~n4892 & ~n5075;
  assign n5077 = n5076 ^ n4884;
  assign n5071 = n4827 ^ n4820;
  assign n5072 = ~n4835 & ~n5071;
  assign n5073 = n5072 ^ n4820;
  assign n5068 = n4907 ^ n4900;
  assign n5069 = ~n4915 & n5068;
  assign n5070 = n5069 ^ n4900;
  assign n5074 = n5073 ^ n5070;
  assign n5078 = n5077 ^ n5074;
  assign n5082 = n5081 ^ n5078;
  assign n5086 = n5085 ^ n5082;
  assign n5090 = n5089 ^ n5086;
  assign n5095 = n5094 ^ n5090;
  assign n5063 = n4852 ^ n4848;
  assign n5064 = ~n4849 & n5063;
  assign n5065 = n5064 ^ n4836;
  assign n5058 = n4874 ^ n4860;
  assign n5059 = n4875 & ~n5058;
  assign n5060 = n5059 ^ n4867;
  assign n5049 = ~x28 & n820;
  assign n5050 = ~x27 & n822;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = x28 & n813;
  assign n5053 = x27 & n817;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = n5051 & n5054;
  assign n5046 = x43 ^ x31;
  assign n5047 = n456 & n5046;
  assign n5048 = ~n460 & ~n5047;
  assign n5056 = n5055 ^ n5048;
  assign n5045 = x10 & x63;
  assign n5057 = n5056 ^ n5045;
  assign n5061 = n5060 ^ n5057;
  assign n5036 = ~x26 & n1037;
  assign n5037 = ~x25 & n1041;
  assign n5038 = ~n5036 & ~n5037;
  assign n5039 = x26 & n1044;
  assign n5040 = x25 & n1046;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n5038 & n5041;
  assign n5029 = ~x18 & n2013;
  assign n5030 = ~x17 & n2017;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = x18 & n2020;
  assign n5033 = x17 & n2022;
  assign n5034 = ~n5032 & ~n5033;
  assign n5035 = n5031 & n5034;
  assign n5043 = n5042 ^ n5035;
  assign n5022 = ~x16 & n2463;
  assign n5023 = ~x15 & n2465;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = x16 & n2456;
  assign n5026 = x15 & n2460;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = n5024 & n5027;
  assign n5044 = n5043 ^ n5028;
  assign n5062 = n5061 ^ n5044;
  assign n5066 = n5065 ^ n5062;
  assign n5017 = n4936 ^ n4927;
  assign n5018 = n4936 ^ n4931;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = n5019 ^ n4927;
  assign n5007 = x24 & n1275;
  assign n5008 = x23 & n1279;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = ~x24 & n1282;
  assign n5011 = ~x23 & n1284;
  assign n5012 = ~n5010 & ~n5011;
  assign n5013 = n5009 & n5012;
  assign n5000 = x14 & n2749;
  assign n5001 = x13 & n2751;
  assign n5002 = ~n5000 & ~n5001;
  assign n5003 = ~x14 & n2742;
  assign n5004 = ~x13 & n2746;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = n5002 & n5005;
  assign n5014 = n5013 ^ n5006;
  assign n4993 = ~x12 & n3163;
  assign n4994 = ~x11 & n3167;
  assign n4995 = ~n4993 & ~n4994;
  assign n4996 = x12 & n3170;
  assign n4997 = x11 & n3172;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n4995 & n4998;
  assign n5015 = n5014 ^ n4999;
  assign n4984 = x22 & n1446;
  assign n4985 = x21 & n1448;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = ~x22 & n1439;
  assign n4988 = ~x21 & n1443;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = n4986 & n4989;
  assign n4977 = ~x20 & n1734;
  assign n4978 = ~x19 & n1738;
  assign n4979 = ~n4977 & ~n4978;
  assign n4980 = x20 & n1741;
  assign n4981 = x19 & n1743;
  assign n4982 = ~n4980 & ~n4981;
  assign n4983 = n4979 & n4982;
  assign n4991 = n4990 ^ n4983;
  assign n4970 = ~x30 & n618;
  assign n4971 = ~x29 & n622;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = x30 & n625;
  assign n4974 = x29 & n627;
  assign n4975 = ~n4973 & ~n4974;
  assign n4976 = n4972 & n4975;
  assign n4992 = n4991 ^ n4976;
  assign n5016 = n5015 ^ n4992;
  assign n5021 = n5020 ^ n5016;
  assign n5067 = n5066 ^ n5021;
  assign n5096 = n5095 ^ n5067;
  assign n5100 = n5099 ^ n5096;
  assign n5104 = n5103 ^ n5100;
  assign n5108 = n5107 ^ n5104;
  assign n5243 = n5107 ^ n5100;
  assign n5244 = ~n5104 & ~n5243;
  assign n5245 = n5244 ^ n5107;
  assign n5239 = n5099 ^ n5095;
  assign n5240 = n5096 & ~n5239;
  assign n5241 = n5240 ^ n5067;
  assign n5235 = n5094 ^ n5089;
  assign n5236 = ~n5090 & n5235;
  assign n5237 = n5236 ^ n5086;
  assign n5229 = n5062 ^ n5021;
  assign n5230 = n5065 ^ n5021;
  assign n5231 = ~n5229 & n5230;
  assign n5232 = n5231 ^ n5062;
  assign n5224 = n5085 ^ n5078;
  assign n5225 = n5085 ^ n5081;
  assign n5226 = ~n5224 & n5225;
  assign n5227 = n5226 ^ n5078;
  assign n5218 = n5077 ^ n5070;
  assign n5219 = n5077 ^ n5073;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = n5220 ^ n5070;
  assign n5214 = n5057 ^ n5044;
  assign n5215 = n5060 ^ n5044;
  assign n5216 = ~n5214 & ~n5215;
  assign n5217 = n5216 ^ n5057;
  assign n5222 = n5221 ^ n5217;
  assign n5210 = n5042 ^ n5028;
  assign n5211 = n5043 & ~n5210;
  assign n5212 = n5211 ^ n5035;
  assign n5206 = n5048 ^ n5045;
  assign n5207 = ~n5056 & ~n5206;
  assign n5208 = n5207 ^ n5045;
  assign n5209 = n5208 ^ n4976;
  assign n5213 = n5212 ^ n5209;
  assign n5223 = n5222 ^ n5213;
  assign n5228 = n5227 ^ n5223;
  assign n5233 = n5232 ^ n5228;
  assign n5202 = n5020 ^ n5015;
  assign n5203 = ~n5016 & n5202;
  assign n5204 = n5203 ^ n4992;
  assign n5196 = n4983 ^ n4976;
  assign n5197 = n4990 ^ n4976;
  assign n5198 = ~n5196 & n5197;
  assign n5199 = n5198 ^ n4983;
  assign n5186 = ~x17 & n2463;
  assign n5187 = ~x16 & n2465;
  assign n5188 = ~n5186 & ~n5187;
  assign n5189 = x17 & n2456;
  assign n5190 = x16 & n2460;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = n5188 & n5191;
  assign n5179 = x19 & n2020;
  assign n5180 = x18 & n2022;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = ~x19 & n2013;
  assign n5183 = ~x18 & n2017;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = n5181 & n5184;
  assign n5193 = n5192 ^ n5185;
  assign n5172 = ~x25 & n1282;
  assign n5173 = ~x24 & n1284;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = x25 & n1275;
  assign n5176 = x24 & n1279;
  assign n5177 = ~n5175 & ~n5176;
  assign n5178 = n5174 & n5177;
  assign n5194 = n5193 ^ n5178;
  assign n5163 = ~x31 & n618;
  assign n5164 = ~x30 & n622;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = x31 & n625;
  assign n5167 = x30 & n627;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = n5165 & n5168;
  assign n5162 = ~n460 & ~n462;
  assign n5170 = n5169 ^ n5162;
  assign n5155 = ~x27 & n1037;
  assign n5156 = ~x26 & n1041;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = x27 & n1044;
  assign n5159 = x26 & n1046;
  assign n5160 = ~n5158 & ~n5159;
  assign n5161 = n5157 & n5160;
  assign n5171 = n5170 ^ n5161;
  assign n5195 = n5194 ^ n5171;
  assign n5200 = n5199 ^ n5195;
  assign n5149 = n5006 ^ n4999;
  assign n5150 = n5013 ^ n4999;
  assign n5151 = n5149 & ~n5150;
  assign n5152 = n5151 ^ n5006;
  assign n5140 = ~x13 & n3163;
  assign n5141 = ~x12 & n3167;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = x13 & n3170;
  assign n5144 = x12 & n3172;
  assign n5145 = ~n5143 & ~n5144;
  assign n5146 = n5142 & n5145;
  assign n5133 = ~x15 & n2742;
  assign n5134 = ~x14 & n2746;
  assign n5135 = ~n5133 & ~n5134;
  assign n5136 = x15 & n2749;
  assign n5137 = x14 & n2751;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = n5135 & n5138;
  assign n5147 = n5146 ^ n5139;
  assign n5126 = ~x29 & n820;
  assign n5127 = ~x28 & n822;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = x29 & n813;
  assign n5130 = x28 & n817;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = n5128 & n5131;
  assign n5148 = n5147 ^ n5132;
  assign n5153 = n5152 ^ n5148;
  assign n5117 = x23 & n1446;
  assign n5118 = x22 & n1448;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = ~x23 & n1439;
  assign n5121 = ~x22 & n1443;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = n5119 & n5122;
  assign n5116 = x11 & x63;
  assign n5124 = n5123 ^ n5116;
  assign n5109 = ~x21 & n1734;
  assign n5110 = ~x20 & n1738;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = x21 & n1741;
  assign n5113 = x20 & n1743;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = n5111 & n5114;
  assign n5125 = n5124 ^ n5115;
  assign n5154 = n5153 ^ n5125;
  assign n5201 = n5200 ^ n5154;
  assign n5205 = n5204 ^ n5201;
  assign n5234 = n5233 ^ n5205;
  assign n5238 = n5237 ^ n5234;
  assign n5242 = n5241 ^ n5238;
  assign n5246 = n5245 ^ n5242;
  assign n5369 = n5245 ^ n5238;
  assign n5370 = n5242 & n5369;
  assign n5371 = n5370 ^ n5245;
  assign n5365 = n5237 ^ n5233;
  assign n5366 = n5234 & ~n5365;
  assign n5367 = n5366 ^ n5205;
  assign n5361 = n5232 ^ n5227;
  assign n5362 = n5228 & n5361;
  assign n5363 = n5362 ^ n5223;
  assign n5356 = n5204 ^ n5200;
  assign n5357 = n5201 & ~n5356;
  assign n5358 = n5357 ^ n5154;
  assign n5352 = n5217 ^ n5213;
  assign n5353 = n5222 & n5352;
  assign n5354 = n5353 ^ n5213;
  assign n5347 = n5212 ^ n5208;
  assign n5348 = ~n5209 & n5347;
  assign n5349 = n5348 ^ n4976;
  assign n5342 = n5139 ^ n5132;
  assign n5343 = n5146 ^ n5132;
  assign n5344 = n5342 & ~n5343;
  assign n5345 = n5344 ^ n5139;
  assign n5334 = ~x20 & n2013;
  assign n5335 = ~x19 & n2017;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = x20 & n2020;
  assign n5338 = x19 & n2022;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = n5336 & n5339;
  assign n5327 = ~x30 & n820;
  assign n5328 = ~x29 & n822;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = x30 & n813;
  assign n5331 = x29 & n817;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = n5329 & n5332;
  assign n5341 = n5340 ^ n5333;
  assign n5346 = n5345 ^ n5341;
  assign n5350 = n5349 ^ n5346;
  assign n5323 = n5192 ^ n5178;
  assign n5324 = n5193 & ~n5323;
  assign n5325 = n5324 ^ n5185;
  assign n5319 = n5169 ^ n5161;
  assign n5320 = ~n5170 & ~n5319;
  assign n5321 = n5320 ^ n5162;
  assign n5316 = n5123 ^ n5115;
  assign n5317 = ~n5124 & ~n5316;
  assign n5318 = n5317 ^ n5116;
  assign n5322 = n5321 ^ n5318;
  assign n5326 = n5325 ^ n5322;
  assign n5351 = n5350 ^ n5326;
  assign n5355 = n5354 ^ n5351;
  assign n5359 = n5358 ^ n5355;
  assign n5311 = n5199 ^ n5194;
  assign n5312 = ~n5195 & ~n5311;
  assign n5313 = n5312 ^ n5171;
  assign n5308 = n5148 ^ n5125;
  assign n5309 = ~n5153 & ~n5308;
  assign n5310 = n5309 ^ n5125;
  assign n5314 = n5313 ^ n5310;
  assign n5297 = x14 & n3170;
  assign n5298 = x13 & n3172;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = ~x14 & n3163;
  assign n5301 = ~x13 & n3167;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = n5299 & n5302;
  assign n5290 = x24 & n1446;
  assign n5291 = x23 & n1448;
  assign n5292 = ~n5290 & ~n5291;
  assign n5293 = ~x24 & n1439;
  assign n5294 = ~x23 & n1443;
  assign n5295 = ~n5293 & ~n5294;
  assign n5296 = n5292 & n5295;
  assign n5304 = n5303 ^ n5296;
  assign n5289 = x12 & x63;
  assign n5305 = n5304 ^ n5289;
  assign n5280 = ~x28 & n1037;
  assign n5281 = ~x27 & n1041;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = x28 & n1044;
  assign n5284 = x27 & n1046;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = n5282 & n5285;
  assign n5277 = x45 ^ x31;
  assign n5278 = n621 & n5277;
  assign n5279 = ~n618 & ~n5278;
  assign n5287 = n5286 ^ n5279;
  assign n5270 = ~x22 & n1734;
  assign n5271 = ~x21 & n1738;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = x22 & n1741;
  assign n5274 = x21 & n1743;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = n5272 & n5275;
  assign n5288 = n5287 ^ n5276;
  assign n5306 = n5305 ^ n5288;
  assign n5261 = x26 & n1275;
  assign n5262 = x25 & n1279;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = ~x26 & n1282;
  assign n5265 = ~x25 & n1284;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n5263 & n5266;
  assign n5254 = x18 & n2456;
  assign n5255 = x17 & n2460;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = ~x18 & n2463;
  assign n5258 = ~x17 & n2465;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = n5256 & n5259;
  assign n5268 = n5267 ^ n5260;
  assign n5247 = ~x16 & n2742;
  assign n5248 = ~x15 & n2746;
  assign n5249 = ~n5247 & ~n5248;
  assign n5250 = x16 & n2749;
  assign n5251 = x15 & n2751;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = n5249 & n5252;
  assign n5269 = n5268 ^ n5253;
  assign n5307 = n5306 ^ n5269;
  assign n5315 = n5314 ^ n5307;
  assign n5360 = n5359 ^ n5315;
  assign n5364 = n5363 ^ n5360;
  assign n5368 = n5367 ^ n5364;
  assign n5372 = n5371 ^ n5368;
  assign n5494 = n5371 ^ n5364;
  assign n5495 = n5368 & ~n5494;
  assign n5496 = n5495 ^ n5371;
  assign n5490 = n5363 ^ n5359;
  assign n5491 = n5360 & n5490;
  assign n5492 = n5491 ^ n5315;
  assign n5486 = n5358 ^ n5354;
  assign n5487 = n5355 & ~n5486;
  assign n5488 = n5487 ^ n5351;
  assign n5482 = n5310 ^ n5307;
  assign n5483 = ~n5314 & n5482;
  assign n5484 = n5483 ^ n5307;
  assign n5476 = n5346 ^ n5326;
  assign n5477 = n5349 ^ n5326;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = n5478 ^ n5346;
  assign n5472 = n5345 ^ n5340;
  assign n5473 = ~n5341 & ~n5472;
  assign n5474 = n5473 ^ n5333;
  assign n5467 = n5325 ^ n5318;
  assign n5468 = n5325 ^ n5321;
  assign n5469 = ~n5467 & n5468;
  assign n5470 = n5469 ^ n5318;
  assign n5458 = x23 & n1741;
  assign n5459 = x22 & n1743;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = ~x23 & n1734;
  assign n5462 = ~x22 & n1738;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = n5460 & n5463;
  assign n5451 = ~x21 & n2013;
  assign n5452 = ~x20 & n2017;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = x21 & n2020;
  assign n5455 = x20 & n2022;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = n5453 & n5456;
  assign n5465 = n5464 ^ n5457;
  assign n5466 = n5465 ^ n5333;
  assign n5471 = n5470 ^ n5466;
  assign n5475 = n5474 ^ n5471;
  assign n5480 = n5479 ^ n5475;
  assign n5445 = n5288 ^ n5269;
  assign n5446 = n5305 ^ n5269;
  assign n5447 = n5445 & n5446;
  assign n5448 = n5447 ^ n5288;
  assign n5441 = n5296 ^ n5289;
  assign n5442 = ~n5304 & ~n5441;
  assign n5443 = n5442 ^ n5289;
  assign n5436 = n5260 ^ n5253;
  assign n5437 = n5267 ^ n5253;
  assign n5438 = n5436 & ~n5437;
  assign n5439 = n5438 ^ n5260;
  assign n5432 = n5279 ^ n5276;
  assign n5433 = n5286 ^ n5276;
  assign n5434 = n5432 & ~n5433;
  assign n5435 = n5434 ^ n5279;
  assign n5440 = n5439 ^ n5435;
  assign n5444 = n5443 ^ n5440;
  assign n5449 = n5448 ^ n5444;
  assign n5421 = x15 & n3170;
  assign n5422 = x14 & n3172;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = ~x15 & n3163;
  assign n5425 = ~x14 & n3167;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = n5423 & n5426;
  assign n5420 = x13 & x63;
  assign n5428 = n5427 ^ n5420;
  assign n5413 = ~x29 & n1037;
  assign n5414 = ~x28 & n1041;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = x29 & n1044;
  assign n5417 = x28 & n1046;
  assign n5418 = ~n5416 & ~n5417;
  assign n5419 = n5415 & n5418;
  assign n5429 = n5428 ^ n5419;
  assign n5404 = ~x17 & n2742;
  assign n5405 = ~x16 & n2746;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = x17 & n2749;
  assign n5408 = x16 & n2751;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = n5406 & n5409;
  assign n5397 = x19 & n2456;
  assign n5398 = x18 & n2460;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = ~x19 & n2463;
  assign n5401 = ~x18 & n2465;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = n5399 & n5402;
  assign n5411 = n5410 ^ n5403;
  assign n5390 = ~x25 & n1439;
  assign n5391 = ~x24 & n1443;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = x25 & n1446;
  assign n5394 = x24 & n1448;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = n5392 & n5395;
  assign n5412 = n5411 ^ n5396;
  assign n5430 = n5429 ^ n5412;
  assign n5381 = ~x31 & n820;
  assign n5382 = ~x30 & n822;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = x31 & n813;
  assign n5385 = x30 & n817;
  assign n5386 = ~n5384 & ~n5385;
  assign n5387 = n5383 & n5386;
  assign n5380 = ~n618 & ~n622;
  assign n5388 = n5387 ^ n5380;
  assign n5373 = x27 & n1275;
  assign n5374 = x26 & n1279;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~x27 & n1282;
  assign n5377 = ~x26 & n1284;
  assign n5378 = ~n5376 & ~n5377;
  assign n5379 = n5375 & n5378;
  assign n5389 = n5388 ^ n5379;
  assign n5431 = n5430 ^ n5389;
  assign n5450 = n5449 ^ n5431;
  assign n5481 = n5480 ^ n5450;
  assign n5485 = n5484 ^ n5481;
  assign n5489 = n5488 ^ n5485;
  assign n5493 = n5492 ^ n5489;
  assign n5497 = n5496 ^ n5493;
  assign n5610 = n5496 ^ n5489;
  assign n5611 = n5493 & ~n5610;
  assign n5612 = n5611 ^ n5496;
  assign n5606 = n5488 ^ n5484;
  assign n5607 = ~n5485 & ~n5606;
  assign n5608 = n5607 ^ n5481;
  assign n5602 = n5475 ^ n5450;
  assign n5603 = n5480 & ~n5602;
  assign n5604 = n5603 ^ n5450;
  assign n5597 = n5448 ^ n5431;
  assign n5598 = n5449 & n5597;
  assign n5599 = n5598 ^ n5431;
  assign n5592 = n5474 ^ n5466;
  assign n5593 = n5474 ^ n5470;
  assign n5594 = ~n5592 & ~n5593;
  assign n5595 = n5594 ^ n5466;
  assign n5588 = n5443 ^ n5439;
  assign n5589 = n5440 & n5588;
  assign n5590 = n5589 ^ n5435;
  assign n5583 = n5457 ^ n5333;
  assign n5584 = n5464 ^ n5333;
  assign n5585 = n5583 & ~n5584;
  assign n5586 = n5585 ^ n5457;
  assign n5574 = ~x28 & n1282;
  assign n5575 = ~x27 & n1284;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = x28 & n1275;
  assign n5578 = x27 & n1279;
  assign n5579 = ~n5577 & ~n5578;
  assign n5580 = n5576 & n5579;
  assign n5567 = ~x22 & n2013;
  assign n5568 = ~x21 & n2017;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = x22 & n2020;
  assign n5571 = x21 & n2022;
  assign n5572 = ~n5570 & ~n5571;
  assign n5573 = n5569 & n5572;
  assign n5581 = n5580 ^ n5573;
  assign n5560 = x20 & n2456;
  assign n5561 = x19 & n2460;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = ~x20 & n2463;
  assign n5564 = ~x19 & n2465;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = n5562 & n5565;
  assign n5582 = n5581 ^ n5566;
  assign n5587 = n5586 ^ n5582;
  assign n5591 = n5590 ^ n5587;
  assign n5596 = n5595 ^ n5591;
  assign n5600 = n5599 ^ n5596;
  assign n5555 = n5412 ^ n5389;
  assign n5556 = n5430 & ~n5555;
  assign n5557 = n5556 ^ n5389;
  assign n5551 = n5403 ^ n5396;
  assign n5552 = ~n5411 & n5551;
  assign n5553 = n5552 ^ n5396;
  assign n5547 = n5387 ^ n5379;
  assign n5548 = ~n5388 & ~n5547;
  assign n5549 = n5548 ^ n5380;
  assign n5544 = x47 ^ x31;
  assign n5545 = n816 & n5544;
  assign n5546 = ~n820 & ~n5545;
  assign n5550 = n5549 ^ n5546;
  assign n5554 = n5553 ^ n5550;
  assign n5558 = n5557 ^ n5554;
  assign n5538 = n5420 ^ n5419;
  assign n5539 = n5427 ^ n5419;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = n5540 ^ n5420;
  assign n5529 = ~x18 & n2742;
  assign n5530 = ~x17 & n2746;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = x18 & n2749;
  assign n5533 = x17 & n2751;
  assign n5534 = ~n5532 & ~n5533;
  assign n5535 = n5531 & n5534;
  assign n5522 = ~x26 & n1439;
  assign n5523 = ~x25 & n1443;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = x26 & n1446;
  assign n5526 = x25 & n1448;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = n5524 & n5527;
  assign n5536 = n5535 ^ n5528;
  assign n5515 = ~x16 & n3163;
  assign n5516 = ~x15 & n3167;
  assign n5517 = ~n5515 & ~n5516;
  assign n5518 = x16 & n3170;
  assign n5519 = x15 & n3172;
  assign n5520 = ~n5518 & ~n5519;
  assign n5521 = n5517 & n5520;
  assign n5537 = n5536 ^ n5521;
  assign n5542 = n5541 ^ n5537;
  assign n5506 = ~x30 & n1037;
  assign n5507 = ~x29 & n1041;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = x30 & n1044;
  assign n5510 = x29 & n1046;
  assign n5511 = ~n5509 & ~n5510;
  assign n5512 = n5508 & n5511;
  assign n5505 = x14 & x63;
  assign n5513 = n5512 ^ n5505;
  assign n5498 = ~x24 & n1734;
  assign n5499 = ~x23 & n1738;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = x24 & n1741;
  assign n5502 = x23 & n1743;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = n5500 & n5503;
  assign n5514 = n5513 ^ n5504;
  assign n5543 = n5542 ^ n5514;
  assign n5559 = n5558 ^ n5543;
  assign n5601 = n5600 ^ n5559;
  assign n5605 = n5604 ^ n5601;
  assign n5609 = n5608 ^ n5605;
  assign n5613 = n5612 ^ n5609;
  assign n5721 = n5612 ^ n5605;
  assign n5722 = ~n5609 & ~n5721;
  assign n5723 = n5722 ^ n5612;
  assign n5717 = n5604 ^ n5600;
  assign n5718 = ~n5601 & n5717;
  assign n5719 = n5718 ^ n5559;
  assign n5712 = n5599 ^ n5591;
  assign n5713 = n5599 ^ n5595;
  assign n5714 = n5712 & ~n5713;
  assign n5715 = n5714 ^ n5591;
  assign n5707 = n5554 ^ n5543;
  assign n5708 = n5558 & n5707;
  assign n5709 = n5708 ^ n5543;
  assign n5703 = n5590 ^ n5586;
  assign n5704 = n5587 & ~n5703;
  assign n5705 = n5704 ^ n5582;
  assign n5698 = n5535 ^ n5521;
  assign n5699 = n5536 & ~n5698;
  assign n5700 = n5699 ^ n5528;
  assign n5690 = x21 & n2456;
  assign n5691 = x20 & n2460;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = ~x21 & n2463;
  assign n5694 = ~x20 & n2465;
  assign n5695 = ~n5693 & ~n5694;
  assign n5696 = n5692 & n5695;
  assign n5697 = n5696 ^ n5546;
  assign n5701 = n5700 ^ n5697;
  assign n5680 = ~x17 & n3163;
  assign n5681 = ~x16 & n3167;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = x17 & n3170;
  assign n5684 = x16 & n3172;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = n5682 & n5685;
  assign n5673 = ~x19 & n2742;
  assign n5674 = ~x18 & n2746;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = x19 & n2749;
  assign n5677 = x18 & n2751;
  assign n5678 = ~n5676 & ~n5677;
  assign n5679 = n5675 & n5678;
  assign n5687 = n5686 ^ n5679;
  assign n5666 = x25 & n1741;
  assign n5667 = x24 & n1743;
  assign n5668 = ~n5666 & ~n5667;
  assign n5669 = ~x25 & n1734;
  assign n5670 = ~x24 & n1738;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = n5668 & n5671;
  assign n5688 = n5687 ^ n5672;
  assign n5657 = ~x31 & n1037;
  assign n5658 = ~x30 & n1041;
  assign n5659 = ~n5657 & ~n5658;
  assign n5660 = x31 & n1044;
  assign n5661 = x30 & n1046;
  assign n5662 = ~n5660 & ~n5661;
  assign n5663 = n5659 & n5662;
  assign n5656 = ~n820 & ~n822;
  assign n5664 = n5663 ^ n5656;
  assign n5649 = ~x27 & n1439;
  assign n5650 = ~x26 & n1443;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = x27 & n1446;
  assign n5653 = x26 & n1448;
  assign n5654 = ~n5652 & ~n5653;
  assign n5655 = n5651 & n5654;
  assign n5665 = n5664 ^ n5655;
  assign n5689 = n5688 ^ n5665;
  assign n5702 = n5701 ^ n5689;
  assign n5706 = n5705 ^ n5702;
  assign n5710 = n5709 ^ n5706;
  assign n5643 = n5553 ^ n5546;
  assign n5644 = n5553 ^ n5549;
  assign n5645 = ~n5643 & n5644;
  assign n5646 = n5645 ^ n5546;
  assign n5640 = n5537 ^ n5514;
  assign n5641 = n5542 & ~n5640;
  assign n5642 = n5641 ^ n5514;
  assign n5647 = n5646 ^ n5642;
  assign n5634 = n5573 ^ n5566;
  assign n5635 = n5580 ^ n5566;
  assign n5636 = n5634 & ~n5635;
  assign n5637 = n5636 ^ n5573;
  assign n5631 = n5512 ^ n5504;
  assign n5632 = ~n5513 & ~n5631;
  assign n5633 = n5632 ^ n5505;
  assign n5638 = n5637 ^ n5633;
  assign n5622 = x29 & n1275;
  assign n5623 = x28 & n1279;
  assign n5624 = ~n5622 & ~n5623;
  assign n5625 = ~x29 & n1282;
  assign n5626 = ~x28 & n1284;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = n5624 & n5627;
  assign n5621 = x15 & x63;
  assign n5629 = n5628 ^ n5621;
  assign n5614 = ~x23 & n2013;
  assign n5615 = ~x22 & n2017;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = x23 & n2020;
  assign n5618 = x22 & n2022;
  assign n5619 = ~n5617 & ~n5618;
  assign n5620 = n5616 & n5619;
  assign n5630 = n5629 ^ n5620;
  assign n5639 = n5638 ^ n5630;
  assign n5648 = n5647 ^ n5639;
  assign n5711 = n5710 ^ n5648;
  assign n5716 = n5715 ^ n5711;
  assign n5720 = n5719 ^ n5716;
  assign n5724 = n5723 ^ n5720;
  assign n5823 = n5723 ^ n5716;
  assign n5824 = ~n5720 & n5823;
  assign n5825 = n5824 ^ n5723;
  assign n5819 = n5715 ^ n5710;
  assign n5820 = ~n5711 & n5819;
  assign n5821 = n5820 ^ n5648;
  assign n5814 = n5709 ^ n5702;
  assign n5815 = n5709 ^ n5705;
  assign n5816 = ~n5814 & ~n5815;
  assign n5817 = n5816 ^ n5702;
  assign n5809 = n5642 ^ n5639;
  assign n5810 = ~n5647 & ~n5809;
  assign n5811 = n5810 ^ n5639;
  assign n5805 = n5701 ^ n5688;
  assign n5806 = ~n5689 & ~n5805;
  assign n5807 = n5806 ^ n5665;
  assign n5794 = x26 & n1741;
  assign n5795 = x25 & n1743;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = ~x26 & n1734;
  assign n5798 = ~x25 & n1738;
  assign n5799 = ~n5797 & ~n5798;
  assign n5800 = n5796 & n5799;
  assign n5787 = ~x18 & n3163;
  assign n5788 = ~x17 & n3167;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = x18 & n3170;
  assign n5791 = x17 & n3172;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = n5789 & n5792;
  assign n5801 = n5800 ^ n5793;
  assign n5786 = x16 & x63;
  assign n5802 = n5801 ^ n5786;
  assign n5777 = x30 & n1275;
  assign n5778 = x29 & n1279;
  assign n5779 = ~n5777 & ~n5778;
  assign n5780 = ~x30 & n1282;
  assign n5781 = ~x29 & n1284;
  assign n5782 = ~n5780 & ~n5781;
  assign n5783 = n5779 & n5782;
  assign n5770 = x24 & n2020;
  assign n5771 = x23 & n2022;
  assign n5772 = ~n5770 & ~n5771;
  assign n5773 = ~x24 & n2013;
  assign n5774 = ~x23 & n2017;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = n5772 & n5775;
  assign n5784 = n5783 ^ n5776;
  assign n5763 = x28 & n1446;
  assign n5764 = x27 & n1448;
  assign n5765 = ~n5763 & ~n5764;
  assign n5766 = ~x28 & n1439;
  assign n5767 = ~x27 & n1443;
  assign n5768 = ~n5766 & ~n5767;
  assign n5769 = n5765 & n5768;
  assign n5785 = n5784 ^ n5769;
  assign n5803 = n5802 ^ n5785;
  assign n5754 = ~x22 & n2463;
  assign n5755 = ~x21 & n2465;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = x22 & n2456;
  assign n5758 = x21 & n2460;
  assign n5759 = ~n5757 & ~n5758;
  assign n5760 = n5756 & n5759;
  assign n5747 = ~x20 & n2742;
  assign n5748 = ~x19 & n2746;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = x20 & n2749;
  assign n5751 = x19 & n2751;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = n5749 & n5752;
  assign n5761 = n5760 ^ n5753;
  assign n5744 = x49 ^ x31;
  assign n5745 = n1040 & n5744;
  assign n5746 = ~n1037 & ~n5745;
  assign n5762 = n5761 ^ n5746;
  assign n5804 = n5803 ^ n5762;
  assign n5808 = n5807 ^ n5804;
  assign n5812 = n5811 ^ n5808;
  assign n5739 = n5633 ^ n5630;
  assign n5740 = n5638 & n5739;
  assign n5741 = n5740 ^ n5630;
  assign n5736 = n5700 ^ n5696;
  assign n5737 = n5697 & ~n5736;
  assign n5738 = n5737 ^ n5546;
  assign n5742 = n5741 ^ n5738;
  assign n5732 = n5628 ^ n5620;
  assign n5733 = ~n5629 & ~n5732;
  assign n5734 = n5733 ^ n5621;
  assign n5728 = n5686 ^ n5672;
  assign n5729 = n5687 & ~n5728;
  assign n5730 = n5729 ^ n5679;
  assign n5725 = n5663 ^ n5655;
  assign n5726 = ~n5664 & ~n5725;
  assign n5727 = n5726 ^ n5656;
  assign n5731 = n5730 ^ n5727;
  assign n5735 = n5734 ^ n5731;
  assign n5743 = n5742 ^ n5735;
  assign n5813 = n5812 ^ n5743;
  assign n5818 = n5817 ^ n5813;
  assign n5822 = n5821 ^ n5818;
  assign n5826 = n5825 ^ n5822;
  assign n5919 = n5825 ^ n5818;
  assign n5920 = n5822 & n5919;
  assign n5921 = n5920 ^ n5825;
  assign n5915 = n5817 ^ n5812;
  assign n5916 = n5813 & ~n5915;
  assign n5917 = n5916 ^ n5743;
  assign n5911 = n5811 ^ n5807;
  assign n5912 = ~n5808 & n5911;
  assign n5913 = n5912 ^ n5804;
  assign n5906 = n5738 ^ n5735;
  assign n5907 = n5742 & n5906;
  assign n5908 = n5907 ^ n5735;
  assign n5902 = n5785 ^ n5762;
  assign n5903 = n5803 & ~n5902;
  assign n5904 = n5903 ^ n5762;
  assign n5891 = ~x31 & n1282;
  assign n5892 = ~x30 & n1284;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = x31 & n1275;
  assign n5895 = x30 & n1279;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = n5893 & n5896;
  assign n5890 = ~n1037 & ~n1041;
  assign n5898 = n5897 ^ n5890;
  assign n5883 = ~x27 & n1734;
  assign n5884 = ~x26 & n1738;
  assign n5885 = ~n5883 & ~n5884;
  assign n5886 = x27 & n1741;
  assign n5887 = x26 & n1743;
  assign n5888 = ~n5886 & ~n5887;
  assign n5889 = n5885 & n5888;
  assign n5899 = n5898 ^ n5889;
  assign n5874 = ~x23 & n2463;
  assign n5875 = ~x22 & n2465;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = x23 & n2456;
  assign n5878 = x22 & n2460;
  assign n5879 = ~n5877 & ~n5878;
  assign n5880 = n5876 & n5879;
  assign n5867 = ~x29 & n1439;
  assign n5868 = ~x28 & n1443;
  assign n5869 = ~n5867 & ~n5868;
  assign n5870 = x29 & n1446;
  assign n5871 = x28 & n1448;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = n5869 & n5872;
  assign n5881 = n5880 ^ n5873;
  assign n5860 = x21 & n2749;
  assign n5861 = x20 & n2751;
  assign n5862 = ~n5860 & ~n5861;
  assign n5863 = ~x21 & n2742;
  assign n5864 = ~x20 & n2746;
  assign n5865 = ~n5863 & ~n5864;
  assign n5866 = n5862 & n5865;
  assign n5882 = n5881 ^ n5866;
  assign n5900 = n5899 ^ n5882;
  assign n5851 = x19 & n3170;
  assign n5852 = x18 & n3172;
  assign n5853 = ~n5851 & ~n5852;
  assign n5854 = ~x19 & n3163;
  assign n5855 = ~x18 & n3167;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = n5853 & n5856;
  assign n5850 = x17 & x63;
  assign n5858 = n5857 ^ n5850;
  assign n5843 = ~x25 & n2013;
  assign n5844 = ~x24 & n2017;
  assign n5845 = ~n5843 & ~n5844;
  assign n5846 = x25 & n2020;
  assign n5847 = x24 & n2022;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = n5845 & n5848;
  assign n5859 = n5858 ^ n5849;
  assign n5901 = n5900 ^ n5859;
  assign n5905 = n5904 ^ n5901;
  assign n5909 = n5908 ^ n5905;
  assign n5838 = n5734 ^ n5727;
  assign n5839 = n5731 & n5838;
  assign n5840 = n5839 ^ n5734;
  assign n5835 = n5753 ^ n5746;
  assign n5836 = ~n5761 & ~n5835;
  assign n5837 = n5836 ^ n5746;
  assign n5841 = n5840 ^ n5837;
  assign n5831 = n5783 ^ n5769;
  assign n5832 = n5784 & ~n5831;
  assign n5833 = n5832 ^ n5776;
  assign n5827 = n5793 ^ n5786;
  assign n5828 = ~n5801 & ~n5827;
  assign n5829 = n5828 ^ n5786;
  assign n5830 = n5829 ^ n5746;
  assign n5834 = n5833 ^ n5830;
  assign n5842 = n5841 ^ n5834;
  assign n5910 = n5909 ^ n5842;
  assign n5914 = n5913 ^ n5910;
  assign n5918 = n5917 ^ n5914;
  assign n5922 = n5921 ^ n5918;
  assign n6011 = n5921 ^ n5914;
  assign n6012 = n5918 & ~n6011;
  assign n6013 = n6012 ^ n5921;
  assign n6007 = n5913 ^ n5909;
  assign n6008 = n5910 & n6007;
  assign n6009 = n6008 ^ n5842;
  assign n6003 = n5908 ^ n5904;
  assign n6004 = ~n5905 & n6003;
  assign n6005 = n6004 ^ n5901;
  assign n5998 = n5837 ^ n5834;
  assign n5999 = n5840 ^ n5834;
  assign n6000 = n5998 & ~n5999;
  assign n6001 = n6000 ^ n5837;
  assign n5993 = n5833 ^ n5829;
  assign n5994 = ~n5830 & n5993;
  assign n5995 = n5994 ^ n5746;
  assign n5987 = n5890 ^ n5889;
  assign n5988 = n5897 ^ n5889;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = n5989 ^ n5890;
  assign n5979 = x20 & n3170;
  assign n5980 = x19 & n3172;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = ~x20 & n3163;
  assign n5983 = ~x19 & n3167;
  assign n5984 = ~n5982 & ~n5983;
  assign n5985 = n5981 & n5984;
  assign n5976 = x51 ^ x31;
  assign n5977 = n1278 & n5976;
  assign n5978 = ~n1282 & ~n5977;
  assign n5986 = n5985 ^ n5978;
  assign n5991 = n5990 ^ n5986;
  assign n5967 = ~x30 & n1439;
  assign n5968 = ~x29 & n1443;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = x30 & n1446;
  assign n5971 = x29 & n1448;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = n5969 & n5972;
  assign n5966 = x18 & x63;
  assign n5974 = n5973 ^ n5966;
  assign n5959 = x26 & n2020;
  assign n5960 = x25 & n2022;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~x26 & n2013;
  assign n5963 = ~x25 & n2017;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = n5961 & n5964;
  assign n5975 = n5974 ^ n5965;
  assign n5992 = n5991 ^ n5975;
  assign n5996 = n5995 ^ n5992;
  assign n5955 = n5899 ^ n5859;
  assign n5956 = ~n5900 & ~n5955;
  assign n5957 = n5956 ^ n5882;
  assign n5950 = n5880 ^ n5866;
  assign n5951 = n5881 & ~n5950;
  assign n5952 = n5951 ^ n5873;
  assign n5946 = n5850 ^ n5849;
  assign n5947 = n5857 ^ n5849;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = n5948 ^ n5850;
  assign n5953 = n5952 ^ n5949;
  assign n5937 = x28 & n1741;
  assign n5938 = x27 & n1743;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = ~x28 & n1734;
  assign n5941 = ~x27 & n1738;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = n5939 & n5942;
  assign n5930 = ~x24 & n2463;
  assign n5931 = ~x23 & n2465;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = x24 & n2456;
  assign n5934 = x23 & n2460;
  assign n5935 = ~n5933 & ~n5934;
  assign n5936 = n5932 & n5935;
  assign n5944 = n5943 ^ n5936;
  assign n5923 = ~x22 & n2742;
  assign n5924 = ~x21 & n2746;
  assign n5925 = ~n5923 & ~n5924;
  assign n5926 = x22 & n2749;
  assign n5927 = x21 & n2751;
  assign n5928 = ~n5926 & ~n5927;
  assign n5929 = n5925 & n5928;
  assign n5945 = n5944 ^ n5929;
  assign n5954 = n5953 ^ n5945;
  assign n5958 = n5957 ^ n5954;
  assign n5997 = n5996 ^ n5958;
  assign n6002 = n6001 ^ n5997;
  assign n6006 = n6005 ^ n6002;
  assign n6010 = n6009 ^ n6006;
  assign n6014 = n6013 ^ n6010;
  assign n6095 = n6013 ^ n6006;
  assign n6096 = ~n6010 & n6095;
  assign n6097 = n6096 ^ n6013;
  assign n6091 = n6005 ^ n6001;
  assign n6092 = ~n6002 & n6091;
  assign n6093 = n6092 ^ n5997;
  assign n6087 = n5996 ^ n5957;
  assign n6088 = ~n5958 & n6087;
  assign n6089 = n6088 ^ n5954;
  assign n6082 = n5995 ^ n5991;
  assign n6083 = ~n5992 & ~n6082;
  assign n6084 = n6083 ^ n5975;
  assign n6078 = n5949 ^ n5945;
  assign n6079 = n5953 & ~n6078;
  assign n6080 = n6079 ^ n5945;
  assign n6073 = n5936 ^ n5929;
  assign n6074 = ~n5944 & n6073;
  assign n6075 = n6074 ^ n5929;
  assign n6070 = n5973 ^ n5965;
  assign n6071 = ~n5974 & ~n6070;
  assign n6072 = n6071 ^ n5966;
  assign n6076 = n6075 ^ n6072;
  assign n6061 = ~x31 & n1439;
  assign n6062 = ~x30 & n1443;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = x31 & n1446;
  assign n6065 = x30 & n1448;
  assign n6066 = ~n6064 & ~n6065;
  assign n6067 = n6063 & n6066;
  assign n6060 = ~n1282 & ~n1284;
  assign n6068 = n6067 ^ n6060;
  assign n6053 = ~x27 & n2013;
  assign n6054 = ~x26 & n2017;
  assign n6055 = ~n6053 & ~n6054;
  assign n6056 = x27 & n2020;
  assign n6057 = x26 & n2022;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = n6055 & n6058;
  assign n6069 = n6068 ^ n6059;
  assign n6077 = n6076 ^ n6069;
  assign n6081 = n6080 ^ n6077;
  assign n6085 = n6084 ^ n6081;
  assign n6049 = n5990 ^ n5985;
  assign n6050 = ~n5986 & n6049;
  assign n6051 = n6050 ^ n5978;
  assign n6039 = ~x25 & n2463;
  assign n6040 = ~x24 & n2465;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = x25 & n2456;
  assign n6043 = x24 & n2460;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = n6041 & n6044;
  assign n6038 = x19 & x63;
  assign n6046 = n6045 ^ n6038;
  assign n6031 = ~x29 & n1734;
  assign n6032 = ~x28 & n1738;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = x29 & n1741;
  assign n6035 = x28 & n1743;
  assign n6036 = ~n6034 & ~n6035;
  assign n6037 = n6033 & n6036;
  assign n6047 = n6046 ^ n6037;
  assign n6022 = ~x21 & n3163;
  assign n6023 = ~x20 & n3167;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = x21 & n3170;
  assign n6026 = x20 & n3172;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = n6024 & n6027;
  assign n6015 = x23 & n2749;
  assign n6016 = x22 & n2751;
  assign n6017 = ~n6015 & ~n6016;
  assign n6018 = ~x23 & n2742;
  assign n6019 = ~x22 & n2746;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n6017 & n6020;
  assign n6029 = n6028 ^ n6021;
  assign n6030 = n6029 ^ n5978;
  assign n6048 = n6047 ^ n6030;
  assign n6052 = n6051 ^ n6048;
  assign n6086 = n6085 ^ n6052;
  assign n6090 = n6089 ^ n6086;
  assign n6094 = n6093 ^ n6090;
  assign n6098 = n6097 ^ n6094;
  assign n6173 = n6097 ^ n6090;
  assign n6174 = ~n6094 & ~n6173;
  assign n6175 = n6174 ^ n6097;
  assign n6168 = n6089 ^ n6052;
  assign n6169 = n6089 ^ n6085;
  assign n6170 = ~n6168 & ~n6169;
  assign n6171 = n6170 ^ n6052;
  assign n6164 = n6084 ^ n6080;
  assign n6165 = n6081 & n6164;
  assign n6166 = n6165 ^ n6077;
  assign n6160 = n6051 ^ n6047;
  assign n6161 = ~n6048 & ~n6160;
  assign n6162 = n6161 ^ n6030;
  assign n6155 = n6072 ^ n6069;
  assign n6156 = n6076 & n6155;
  assign n6157 = n6156 ^ n6069;
  assign n6151 = n6045 ^ n6037;
  assign n6152 = ~n6046 & ~n6151;
  assign n6153 = n6152 ^ n6038;
  assign n6147 = n6067 ^ n6059;
  assign n6148 = ~n6068 & ~n6147;
  assign n6149 = n6148 ^ n6060;
  assign n6144 = x53 ^ x31;
  assign n6145 = n1442 & n6144;
  assign n6146 = ~n1439 & ~n6145;
  assign n6150 = n6149 ^ n6146;
  assign n6154 = n6153 ^ n6150;
  assign n6158 = n6157 ^ n6154;
  assign n6140 = n6021 ^ n5978;
  assign n6141 = ~n6029 & n6140;
  assign n6142 = n6141 ^ n5978;
  assign n6130 = x26 & n2456;
  assign n6131 = x25 & n2460;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = ~x26 & n2463;
  assign n6134 = ~x25 & n2465;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = n6132 & n6135;
  assign n6123 = ~x30 & n1734;
  assign n6124 = ~x29 & n1738;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = x30 & n1741;
  assign n6127 = x29 & n1743;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = n6125 & n6128;
  assign n6137 = n6136 ^ n6129;
  assign n6116 = ~x24 & n2742;
  assign n6117 = ~x23 & n2746;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = x24 & n2749;
  assign n6120 = x23 & n2751;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = n6118 & n6121;
  assign n6138 = n6137 ^ n6122;
  assign n6107 = ~x22 & n3163;
  assign n6108 = ~x21 & n3167;
  assign n6109 = ~n6107 & ~n6108;
  assign n6110 = x22 & n3170;
  assign n6111 = x21 & n3172;
  assign n6112 = ~n6110 & ~n6111;
  assign n6113 = n6109 & n6112;
  assign n6100 = ~x28 & n2013;
  assign n6101 = ~x27 & n2017;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = x28 & n2020;
  assign n6104 = x27 & n2022;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = n6102 & n6105;
  assign n6114 = n6113 ^ n6106;
  assign n6099 = x20 & x63;
  assign n6115 = n6114 ^ n6099;
  assign n6139 = n6138 ^ n6115;
  assign n6143 = n6142 ^ n6139;
  assign n6159 = n6158 ^ n6143;
  assign n6163 = n6162 ^ n6159;
  assign n6167 = n6166 ^ n6163;
  assign n6172 = n6171 ^ n6167;
  assign n6176 = n6175 ^ n6172;
  assign n6246 = n6175 ^ n6167;
  assign n6247 = n6172 & n6246;
  assign n6248 = n6247 ^ n6175;
  assign n6242 = n6166 ^ n6162;
  assign n6243 = ~n6163 & ~n6242;
  assign n6244 = n6243 ^ n6159;
  assign n6238 = n6154 ^ n6143;
  assign n6239 = ~n6158 & n6238;
  assign n6240 = n6239 ^ n6143;
  assign n6233 = n6142 ^ n6138;
  assign n6234 = ~n6139 & ~n6233;
  assign n6235 = n6234 ^ n6115;
  assign n6228 = n6153 ^ n6146;
  assign n6229 = n6153 ^ n6149;
  assign n6230 = n6228 & ~n6229;
  assign n6231 = n6230 ^ n6146;
  assign n6224 = n6136 ^ n6122;
  assign n6225 = n6137 & ~n6224;
  assign n6226 = n6225 ^ n6129;
  assign n6222 = x21 & x63;
  assign n6223 = n6222 ^ n6146;
  assign n6227 = n6226 ^ n6223;
  assign n6232 = n6231 ^ n6227;
  assign n6236 = n6235 ^ n6232;
  assign n6217 = n6106 ^ n6099;
  assign n6218 = ~n6114 & ~n6217;
  assign n6219 = n6218 ^ n6099;
  assign n6208 = x29 & n2020;
  assign n6209 = x28 & n2022;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = ~x29 & n2013;
  assign n6212 = ~x28 & n2017;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = n6210 & n6213;
  assign n6201 = ~x25 & n2742;
  assign n6202 = ~x24 & n2746;
  assign n6203 = ~n6201 & ~n6202;
  assign n6204 = x25 & n2749;
  assign n6205 = x24 & n2751;
  assign n6206 = ~n6204 & ~n6205;
  assign n6207 = n6203 & n6206;
  assign n6215 = n6214 ^ n6207;
  assign n6194 = x23 & n3170;
  assign n6195 = x22 & n3172;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = ~x23 & n3163;
  assign n6198 = ~x22 & n3167;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = n6196 & n6199;
  assign n6216 = n6215 ^ n6200;
  assign n6220 = n6219 ^ n6216;
  assign n6185 = x31 & n1741;
  assign n6186 = x30 & n1743;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = ~x31 & n1734;
  assign n6189 = ~x30 & n1738;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = n6187 & n6190;
  assign n6184 = ~n1439 & ~n1443;
  assign n6192 = n6191 ^ n6184;
  assign n6177 = ~x27 & n2463;
  assign n6178 = ~x26 & n2465;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = x27 & n2456;
  assign n6181 = x26 & n2460;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = n6179 & n6182;
  assign n6193 = n6192 ^ n6183;
  assign n6221 = n6220 ^ n6193;
  assign n6237 = n6236 ^ n6221;
  assign n6241 = n6240 ^ n6237;
  assign n6245 = n6244 ^ n6241;
  assign n6249 = n6248 ^ n6245;
  assign n6314 = n6248 ^ n6241;
  assign n6315 = n6245 & ~n6314;
  assign n6316 = n6315 ^ n6248;
  assign n6310 = n6240 ^ n6236;
  assign n6311 = ~n6237 & ~n6310;
  assign n6312 = n6311 ^ n6221;
  assign n6305 = n6235 ^ n6227;
  assign n6306 = n6235 ^ n6231;
  assign n6307 = n6305 & ~n6306;
  assign n6308 = n6307 ^ n6227;
  assign n6299 = n6216 ^ n6193;
  assign n6300 = n6219 ^ n6193;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = n6301 ^ n6216;
  assign n6295 = n6226 ^ n6146;
  assign n6296 = ~n6223 & ~n6295;
  assign n6297 = n6296 ^ n6222;
  assign n6286 = ~x28 & n2463;
  assign n6287 = ~x27 & n2465;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = x28 & n2456;
  assign n6290 = x27 & n2460;
  assign n6291 = ~n6289 & ~n6290;
  assign n6292 = n6288 & n6291;
  assign n6285 = x22 & x63;
  assign n6293 = n6292 ^ n6285;
  assign n6278 = x30 & n2020;
  assign n6279 = x29 & n2022;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = ~x30 & n2013;
  assign n6282 = ~x29 & n2017;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = n6280 & n6283;
  assign n6294 = n6293 ^ n6284;
  assign n6298 = n6297 ^ n6294;
  assign n6303 = n6302 ^ n6298;
  assign n6272 = n6207 ^ n6200;
  assign n6273 = n6214 ^ n6200;
  assign n6274 = n6272 & ~n6273;
  assign n6275 = n6274 ^ n6207;
  assign n6269 = n6191 ^ n6183;
  assign n6270 = ~n6192 & ~n6269;
  assign n6271 = n6270 ^ n6184;
  assign n6276 = n6275 ^ n6271;
  assign n6260 = ~x26 & n2742;
  assign n6261 = ~x25 & n2746;
  assign n6262 = ~n6260 & ~n6261;
  assign n6263 = x26 & n2749;
  assign n6264 = x25 & n2751;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = n6262 & n6265;
  assign n6253 = x24 & n3170;
  assign n6254 = x23 & n3172;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~x24 & n3163;
  assign n6257 = ~x23 & n3167;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259 = n6255 & n6258;
  assign n6267 = n6266 ^ n6259;
  assign n6250 = x55 ^ x31;
  assign n6251 = n1737 & n6250;
  assign n6252 = ~n1734 & ~n6251;
  assign n6268 = n6267 ^ n6252;
  assign n6277 = n6276 ^ n6268;
  assign n6304 = n6303 ^ n6277;
  assign n6309 = n6308 ^ n6304;
  assign n6313 = n6312 ^ n6309;
  assign n6317 = n6316 ^ n6313;
  assign n6375 = n6316 ^ n6309;
  assign n6376 = n6313 & n6375;
  assign n6377 = n6376 ^ n6316;
  assign n6371 = n6308 ^ n6303;
  assign n6372 = n6304 & ~n6371;
  assign n6373 = n6372 ^ n6277;
  assign n6367 = n6302 ^ n6297;
  assign n6368 = ~n6298 & n6367;
  assign n6369 = n6368 ^ n6294;
  assign n6363 = n6271 ^ n6268;
  assign n6364 = n6276 & ~n6363;
  assign n6365 = n6364 ^ n6268;
  assign n6357 = n6285 ^ n6284;
  assign n6358 = n6292 ^ n6284;
  assign n6359 = n6357 & n6358;
  assign n6360 = n6359 ^ n6285;
  assign n6348 = ~x31 & n2013;
  assign n6349 = ~x30 & n2017;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = x31 & n2020;
  assign n6352 = x30 & n2022;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = n6350 & n6353;
  assign n6347 = ~n1734 & ~n1738;
  assign n6355 = n6354 ^ n6347;
  assign n6340 = ~x27 & n2742;
  assign n6341 = ~x26 & n2746;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = x27 & n2749;
  assign n6344 = x26 & n2751;
  assign n6345 = ~n6343 & ~n6344;
  assign n6346 = n6342 & n6345;
  assign n6356 = n6355 ^ n6346;
  assign n6361 = n6360 ^ n6356;
  assign n6335 = n6259 ^ n6252;
  assign n6336 = ~n6267 & n6335;
  assign n6337 = n6336 ^ n6252;
  assign n6338 = n6337 ^ n6284;
  assign n6326 = ~x25 & n3163;
  assign n6327 = ~x24 & n3167;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = x25 & n3170;
  assign n6330 = x24 & n3172;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = n6328 & n6331;
  assign n6319 = x29 & n2456;
  assign n6320 = x28 & n2460;
  assign n6321 = ~n6319 & ~n6320;
  assign n6322 = ~x29 & n2463;
  assign n6323 = ~x28 & n2465;
  assign n6324 = ~n6322 & ~n6323;
  assign n6325 = n6321 & n6324;
  assign n6333 = n6332 ^ n6325;
  assign n6318 = x23 & x63;
  assign n6334 = n6333 ^ n6318;
  assign n6339 = n6338 ^ n6334;
  assign n6362 = n6361 ^ n6339;
  assign n6366 = n6365 ^ n6362;
  assign n6370 = n6369 ^ n6366;
  assign n6374 = n6373 ^ n6370;
  assign n6378 = n6377 ^ n6374;
  assign n6429 = n6377 ^ n6370;
  assign n6430 = ~n6374 & n6429;
  assign n6431 = n6430 ^ n6377;
  assign n6425 = n6369 ^ n6365;
  assign n6426 = ~n6366 & ~n6425;
  assign n6427 = n6426 ^ n6362;
  assign n6421 = n6360 ^ n6339;
  assign n6422 = n6361 & ~n6421;
  assign n6423 = n6422 ^ n6356;
  assign n6416 = n6334 ^ n6284;
  assign n6417 = n6337 ^ n6334;
  assign n6418 = ~n6416 & n6417;
  assign n6419 = n6418 ^ n6284;
  assign n6411 = n6354 ^ n6346;
  assign n6412 = ~n6355 & ~n6411;
  assign n6413 = n6412 ^ n6347;
  assign n6402 = x26 & n3170;
  assign n6403 = x25 & n3172;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~x26 & n3163;
  assign n6406 = ~x25 & n3167;
  assign n6407 = ~n6405 & ~n6406;
  assign n6408 = n6404 & n6407;
  assign n6401 = x24 & x63;
  assign n6409 = n6408 ^ n6401;
  assign n6398 = x57 ^ x31;
  assign n6399 = n2016 & n6398;
  assign n6400 = ~n2013 & ~n6399;
  assign n6410 = n6409 ^ n6400;
  assign n6414 = n6413 ^ n6410;
  assign n6394 = n6325 ^ n6318;
  assign n6395 = ~n6333 & ~n6394;
  assign n6396 = n6395 ^ n6318;
  assign n6386 = ~x28 & n2742;
  assign n6387 = ~x27 & n2746;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = x28 & n2749;
  assign n6390 = x27 & n2751;
  assign n6391 = ~n6389 & ~n6390;
  assign n6392 = n6388 & n6391;
  assign n6379 = ~x30 & n2463;
  assign n6380 = ~x29 & n2465;
  assign n6381 = ~n6379 & ~n6380;
  assign n6382 = x30 & n2456;
  assign n6383 = x29 & n2460;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = n6381 & n6384;
  assign n6393 = n6392 ^ n6385;
  assign n6397 = n6396 ^ n6393;
  assign n6415 = n6414 ^ n6397;
  assign n6420 = n6419 ^ n6415;
  assign n6424 = n6423 ^ n6420;
  assign n6428 = n6427 ^ n6424;
  assign n6432 = n6431 ^ n6428;
  assign n6478 = n6431 ^ n6424;
  assign n6479 = ~n6428 & n6478;
  assign n6480 = n6479 ^ n6431;
  assign n6474 = n6423 ^ n6419;
  assign n6475 = n6420 & n6474;
  assign n6476 = n6475 ^ n6415;
  assign n6470 = n6413 ^ n6397;
  assign n6471 = n6414 & n6470;
  assign n6472 = n6471 ^ n6410;
  assign n6466 = n6396 ^ n6392;
  assign n6467 = ~n6393 & n6466;
  assign n6468 = n6467 ^ n6385;
  assign n6460 = n6401 ^ n6400;
  assign n6461 = n6408 ^ n6400;
  assign n6462 = ~n6460 & ~n6461;
  assign n6463 = n6462 ^ n6401;
  assign n6451 = ~x31 & n2463;
  assign n6452 = ~x30 & n2465;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = x31 & n2456;
  assign n6455 = x30 & n2460;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = n6453 & n6456;
  assign n6450 = ~n2013 & ~n2017;
  assign n6458 = n6457 ^ n6450;
  assign n6443 = x27 & n3170;
  assign n6444 = x26 & n3172;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = ~x27 & n3163;
  assign n6447 = ~x26 & n3167;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = n6445 & n6448;
  assign n6459 = n6458 ^ n6449;
  assign n6464 = n6463 ^ n6459;
  assign n6434 = ~x29 & n2742;
  assign n6435 = ~x28 & n2746;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = x29 & n2749;
  assign n6438 = x28 & n2751;
  assign n6439 = ~n6437 & ~n6438;
  assign n6440 = n6436 & n6439;
  assign n6433 = x25 & x63;
  assign n6441 = n6440 ^ n6433;
  assign n6442 = n6441 ^ n6385;
  assign n6465 = n6464 ^ n6442;
  assign n6469 = n6468 ^ n6465;
  assign n6473 = n6472 ^ n6469;
  assign n6477 = n6476 ^ n6473;
  assign n6481 = n6480 ^ n6477;
  assign n6521 = n6480 ^ n6473;
  assign n6522 = n6477 & n6521;
  assign n6523 = n6522 ^ n6480;
  assign n6517 = n6472 ^ n6468;
  assign n6518 = n6469 & ~n6517;
  assign n6519 = n6518 ^ n6465;
  assign n6513 = n6459 ^ n6442;
  assign n6514 = ~n6464 & n6513;
  assign n6515 = n6514 ^ n6442;
  assign n6508 = n6433 ^ n6385;
  assign n6509 = n6440 ^ n6385;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = n6510 ^ n6433;
  assign n6502 = n6450 ^ n6449;
  assign n6503 = n6457 ^ n6449;
  assign n6504 = ~n6502 & ~n6503;
  assign n6505 = n6504 ^ n6450;
  assign n6499 = x59 ^ x31;
  assign n6500 = n2459 & n6499;
  assign n6501 = ~n2463 & ~n6500;
  assign n6506 = n6505 ^ n6501;
  assign n6490 = ~x30 & n2742;
  assign n6491 = ~x29 & n2746;
  assign n6492 = ~n6490 & ~n6491;
  assign n6493 = x30 & n2749;
  assign n6494 = x29 & n2751;
  assign n6495 = ~n6493 & ~n6494;
  assign n6496 = n6492 & n6495;
  assign n6489 = x26 & x63;
  assign n6497 = n6496 ^ n6489;
  assign n6482 = x28 & n3170;
  assign n6483 = x27 & n3172;
  assign n6484 = ~n6482 & ~n6483;
  assign n6485 = ~x28 & n3163;
  assign n6486 = ~x27 & n3167;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = n6484 & n6487;
  assign n6498 = n6497 ^ n6488;
  assign n6507 = n6506 ^ n6498;
  assign n6512 = n6511 ^ n6507;
  assign n6516 = n6515 ^ n6512;
  assign n6520 = n6519 ^ n6516;
  assign n6524 = n6523 ^ n6520;
  assign n6558 = n6523 ^ n6516;
  assign n6559 = ~n6520 & n6558;
  assign n6560 = n6559 ^ n6523;
  assign n6554 = n6515 ^ n6507;
  assign n6555 = n6512 & ~n6554;
  assign n6556 = n6555 ^ n6511;
  assign n6549 = n6501 ^ n6498;
  assign n6550 = n6505 ^ n6498;
  assign n6551 = n6549 & ~n6550;
  assign n6552 = n6551 ^ n6501;
  assign n6544 = n6496 ^ n6488;
  assign n6545 = ~n6497 & ~n6544;
  assign n6546 = n6545 ^ n6489;
  assign n6536 = ~x29 & n3163;
  assign n6537 = ~x28 & n3167;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = x29 & n3170;
  assign n6540 = x28 & n3172;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = n6538 & n6541;
  assign n6543 = n6542 ^ n6501;
  assign n6547 = n6546 ^ n6543;
  assign n6527 = x31 & n2749;
  assign n6528 = x30 & n2751;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = ~x31 & n2742;
  assign n6531 = ~x30 & n2746;
  assign n6532 = ~n6530 & ~n6531;
  assign n6533 = n6529 & n6532;
  assign n6526 = ~n2463 & ~n2465;
  assign n6534 = n6533 ^ n6526;
  assign n6525 = x27 & x63;
  assign n6535 = n6534 ^ n6525;
  assign n6548 = n6547 ^ n6535;
  assign n6553 = n6552 ^ n6548;
  assign n6557 = n6556 ^ n6553;
  assign n6561 = n6560 ^ n6557;
  assign n6587 = n6560 ^ n6553;
  assign n6588 = n6557 & ~n6587;
  assign n6589 = n6588 ^ n6560;
  assign n6583 = n6552 ^ n6547;
  assign n6584 = ~n6548 & ~n6583;
  assign n6585 = n6584 ^ n6535;
  assign n6579 = n6546 ^ n6542;
  assign n6580 = n6543 & n6579;
  assign n6581 = n6580 ^ n6501;
  assign n6575 = n6526 ^ n6525;
  assign n6576 = n6534 & n6575;
  assign n6577 = n6576 ^ n6525;
  assign n6566 = ~x30 & n3163;
  assign n6567 = ~x29 & n3167;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = x30 & n3170;
  assign n6570 = x29 & n3172;
  assign n6571 = ~n6569 & ~n6570;
  assign n6572 = n6568 & n6571;
  assign n6565 = x28 & x63;
  assign n6573 = n6572 ^ n6565;
  assign n6562 = x61 ^ x31;
  assign n6563 = n2745 & n6562;
  assign n6564 = ~n2742 & ~n6563;
  assign n6574 = n6573 ^ n6564;
  assign n6578 = n6577 ^ n6574;
  assign n6582 = n6581 ^ n6578;
  assign n6586 = n6585 ^ n6582;
  assign n6590 = n6589 ^ n6586;
  assign n6612 = n6589 ^ n6582;
  assign n6613 = n6586 & n6612;
  assign n6614 = n6613 ^ n6589;
  assign n6608 = n6581 ^ n6577;
  assign n6609 = ~n6578 & n6608;
  assign n6610 = n6609 ^ n6574;
  assign n6603 = n6565 ^ n6564;
  assign n6604 = n6572 ^ n6564;
  assign n6605 = n6603 & n6604;
  assign n6606 = n6605 ^ n6565;
  assign n6593 = x31 & n3170;
  assign n6594 = x30 & n3172;
  assign n6595 = ~n6593 & ~n6594;
  assign n6596 = ~x31 & n3163;
  assign n6597 = ~x30 & n3167;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = n6595 & n6598;
  assign n6592 = ~n2742 & ~n2746;
  assign n6600 = n6599 ^ n6592;
  assign n6591 = x29 & x63;
  assign n6601 = n6600 ^ n6591;
  assign n6602 = n6601 ^ n6564;
  assign n6607 = n6606 ^ n6602;
  assign n6611 = n6610 ^ n6607;
  assign n6615 = n6614 ^ n6611;
  assign n6629 = n6614 ^ n6607;
  assign n6630 = n6611 & n6629;
  assign n6631 = n6630 ^ n6614;
  assign n6625 = n6606 ^ n6601;
  assign n6626 = n6602 & n6625;
  assign n6627 = n6626 ^ n6564;
  assign n6621 = n6592 ^ n6591;
  assign n6622 = n6600 & n6621;
  assign n6623 = n6622 ^ n6591;
  assign n6617 = x63 ^ x31;
  assign n6618 = n3166 & n6617;
  assign n6619 = ~n3163 & ~n6618;
  assign n6616 = x30 & x63;
  assign n6620 = n6619 ^ n6616;
  assign n6624 = n6623 ^ n6620;
  assign n6628 = n6627 ^ n6624;
  assign n6632 = n6631 ^ n6628;
  assign n6641 = n6631 ^ n6624;
  assign n6642 = n6628 & n6641;
  assign n6643 = n6642 ^ n6631;
  assign n6637 = n6623 ^ n6619;
  assign n6638 = n6620 & n6637;
  assign n6639 = n6638 ^ n6616;
  assign n6633 = ~n2887 & ~n3166;
  assign n6634 = n6633 ^ x31;
  assign n6635 = x63 & ~n6634;
  assign n6636 = n6635 ^ n6616;
  assign n6640 = n6639 ^ n6636;
  assign n6644 = n6643 ^ n6640;
  assign y0 = n65;
  assign y1 = ~n77;
  assign y2 = ~n88;
  assign y3 = n117;
  assign y4 = n140;
  assign y5 = ~n182;
  assign y6 = n217;
  assign y7 = ~n270;
  assign y8 = n319;
  assign y9 = n385;
  assign y10 = n445;
  assign y11 = n523;
  assign y12 = n594;
  assign y13 = ~n684;
  assign y14 = ~n767;
  assign y15 = ~n869;
  assign y16 = ~n967;
  assign y17 = ~n1081;
  assign y18 = n1189;
  assign y19 = n1315;
  assign y20 = ~n1438;
  assign y21 = n1577;
  assign y22 = ~n1710;
  assign y23 = ~n1861;
  assign y24 = ~n2005;
  assign y25 = n2170;
  assign y26 = ~n2329;
  assign y27 = n2505;
  assign y28 = n2675;
  assign y29 = n2863;
  assign y30 = n3044;
  assign y31 = ~n3244;
  assign y32 = n3431;
  assign y33 = ~n3621;
  assign y34 = n3807;
  assign y35 = ~n3991;
  assign y36 = ~n4171;
  assign y37 = n4345;
  assign y38 = ~n4508;
  assign y39 = ~n4667;
  assign y40 = ~n4819;
  assign y41 = n4969;
  assign y42 = n5108;
  assign y43 = ~n5246;
  assign y44 = ~n5372;
  assign y45 = ~n5497;
  assign y46 = n5613;
  assign y47 = n5724;
  assign y48 = ~n5826;
  assign y49 = ~n5922;
  assign y50 = n6014;
  assign y51 = n6098;
  assign y52 = ~n6176;
  assign y53 = ~n6249;
  assign y54 = ~n6317;
  assign y55 = n6378;
  assign y56 = n6432;
  assign y57 = ~n6481;
  assign y58 = n6524;
  assign y59 = ~n6561;
  assign y60 = ~n6590;
  assign y61 = ~n6615;
  assign y62 = ~n6632;
  assign y63 = n6644;
endmodule