module Xor(
    //output logic out
);

    logic a;
    logic b;

    assign a = 0;
    assign b = 1;

    //assign out = a ^ b;
    
endmodule
