module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288;
  assign n65 = ~x29 & x61;
  assign n66 = ~x28 & x60;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~x30 & x62;
  assign n69 = ~x31 & x63;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & n70;
  assign n72 = ~x25 & x57;
  assign n73 = ~x26 & x58;
  assign n74 = ~x27 & x59;
  assign n75 = ~n73 & ~n74;
  assign n76 = ~n72 & n75;
  assign n77 = ~x56 & n76;
  assign n78 = x24 & n77;
  assign n79 = x59 ^ x27;
  assign n80 = x58 ^ x26;
  assign n81 = n80 ^ n74;
  assign n82 = x57 ^ x25;
  assign n83 = ~x57 & ~n82;
  assign n84 = n83 ^ x26;
  assign n85 = n84 ^ x57;
  assign n86 = n81 & ~n85;
  assign n87 = n86 ^ n83;
  assign n88 = n87 ^ x57;
  assign n89 = n88 ^ x59;
  assign n90 = ~n79 & n89;
  assign n91 = n90 ^ x59;
  assign n92 = ~n78 & n91;
  assign n93 = n71 & ~n92;
  assign n94 = x24 & n76;
  assign n95 = ~n77 & ~n94;
  assign n96 = n71 & ~n95;
  assign n97 = ~x22 & x54;
  assign n98 = ~x23 & x55;
  assign n99 = ~n97 & ~n98;
  assign n100 = x53 ^ x21;
  assign n101 = x53 ^ x20;
  assign n102 = n101 ^ x53;
  assign n103 = x53 ^ x52;
  assign n104 = n103 ^ x53;
  assign n105 = n102 & ~n104;
  assign n106 = n105 ^ x53;
  assign n107 = ~n100 & n106;
  assign n108 = n107 ^ x21;
  assign n109 = n99 & n108;
  assign n110 = ~x21 & x53;
  assign n111 = ~x20 & x52;
  assign n112 = ~n110 & ~n111;
  assign n113 = n99 & n112;
  assign n114 = x51 ^ x19;
  assign n115 = x49 ^ x17;
  assign n116 = x49 ^ x16;
  assign n117 = n116 ^ x49;
  assign n118 = x49 ^ x48;
  assign n119 = n118 ^ x49;
  assign n120 = n117 & ~n119;
  assign n121 = n120 ^ x49;
  assign n122 = ~n115 & n121;
  assign n123 = n122 ^ x17;
  assign n124 = n123 ^ x51;
  assign n125 = n124 ^ x51;
  assign n126 = ~x18 & x50;
  assign n127 = n126 ^ x51;
  assign n128 = n127 ^ x51;
  assign n129 = n125 & ~n128;
  assign n130 = n129 ^ x51;
  assign n133 = n130 ^ x51;
  assign n131 = n130 ^ x50;
  assign n132 = n131 ^ n130;
  assign n134 = n133 ^ n132;
  assign n135 = n130 ^ x18;
  assign n136 = n135 ^ n130;
  assign n137 = n136 ^ n132;
  assign n138 = ~n132 & ~n137;
  assign n139 = n138 ^ n132;
  assign n140 = n134 & ~n139;
  assign n141 = n140 ^ n138;
  assign n142 = n141 ^ n130;
  assign n143 = n142 ^ n132;
  assign n144 = ~n114 & ~n143;
  assign n145 = n144 ^ x19;
  assign n146 = n113 & n145;
  assign n147 = ~n109 & ~n146;
  assign n148 = x55 ^ x23;
  assign n149 = x55 ^ x22;
  assign n150 = n149 ^ x55;
  assign n151 = x55 ^ x54;
  assign n152 = n151 ^ x55;
  assign n153 = n150 & ~n152;
  assign n154 = n153 ^ x55;
  assign n155 = ~n148 & n154;
  assign n156 = n155 ^ x23;
  assign n157 = n147 & ~n156;
  assign n158 = n96 & ~n157;
  assign n159 = ~n93 & ~n158;
  assign n160 = ~x17 & x49;
  assign n161 = ~x19 & x51;
  assign n162 = ~n126 & ~n161;
  assign n163 = ~x16 & x48;
  assign n164 = ~x13 & x45;
  assign n165 = ~x15 & x47;
  assign n166 = ~x14 & x46;
  assign n167 = ~n165 & ~n166;
  assign n168 = ~n164 & n167;
  assign n169 = ~x12 & x44;
  assign n170 = ~x11 & x43;
  assign n171 = ~x10 & x42;
  assign n172 = ~n170 & ~n171;
  assign n173 = ~x9 & x41;
  assign n174 = ~x40 & ~n173;
  assign n175 = n172 & n174;
  assign n176 = x8 & ~n173;
  assign n177 = n172 & n176;
  assign n178 = ~n175 & ~n177;
  assign n179 = x39 ^ x7;
  assign n180 = x39 ^ x6;
  assign n181 = n180 ^ x39;
  assign n182 = x39 ^ x38;
  assign n183 = n182 ^ x39;
  assign n184 = n181 & ~n183;
  assign n185 = n184 ^ x39;
  assign n186 = ~n179 & n185;
  assign n187 = n186 ^ x7;
  assign n188 = ~x6 & x38;
  assign n189 = ~x7 & x39;
  assign n190 = ~n188 & ~n189;
  assign n191 = x37 ^ x5;
  assign n192 = x36 ^ x4;
  assign n193 = x35 ^ x3;
  assign n194 = x34 ^ x2;
  assign n196 = ~x2 & x34;
  assign n195 = x33 ^ x1;
  assign n197 = n196 ^ n195;
  assign n198 = x32 ^ x0;
  assign n199 = x32 & ~n198;
  assign n200 = n199 ^ x1;
  assign n201 = n200 ^ x32;
  assign n202 = n197 & ~n201;
  assign n203 = n202 ^ n199;
  assign n204 = n203 ^ x32;
  assign n205 = n204 ^ x34;
  assign n206 = ~n194 & n205;
  assign n207 = n206 ^ x34;
  assign n208 = n207 ^ x35;
  assign n209 = ~n193 & n208;
  assign n210 = n209 ^ x35;
  assign n211 = n210 ^ x36;
  assign n212 = ~n192 & n211;
  assign n213 = n212 ^ x36;
  assign n214 = n213 ^ x37;
  assign n215 = ~n191 & n214;
  assign n216 = n215 ^ x37;
  assign n217 = n190 & ~n216;
  assign n218 = ~n187 & ~n217;
  assign n219 = ~n178 & ~n218;
  assign n220 = x8 & n175;
  assign n221 = x43 ^ x11;
  assign n222 = x42 ^ x10;
  assign n223 = x9 & ~x41;
  assign n224 = n223 ^ x42;
  assign n225 = ~n222 & ~n224;
  assign n226 = n225 ^ x42;
  assign n227 = n226 ^ x43;
  assign n228 = ~n221 & n227;
  assign n229 = n228 ^ x43;
  assign n230 = ~n220 & n229;
  assign n231 = ~n219 & n230;
  assign n232 = ~n169 & ~n231;
  assign n233 = n168 & n232;
  assign n234 = x12 & n168;
  assign n235 = ~x44 & n234;
  assign n236 = x47 ^ x15;
  assign n237 = x46 ^ x14;
  assign n238 = n237 ^ n165;
  assign n239 = x45 ^ x13;
  assign n240 = ~x45 & ~n239;
  assign n241 = n240 ^ x14;
  assign n242 = n241 ^ x45;
  assign n243 = n238 & ~n242;
  assign n244 = n243 ^ n240;
  assign n245 = n244 ^ x45;
  assign n246 = n245 ^ x47;
  assign n247 = ~n236 & n246;
  assign n248 = n247 ^ x47;
  assign n249 = ~n235 & n248;
  assign n250 = ~n233 & n249;
  assign n251 = ~n163 & ~n250;
  assign n252 = n162 & n251;
  assign n253 = ~n160 & n252;
  assign n254 = n113 & n253;
  assign n255 = n96 & n254;
  assign n256 = x63 ^ x31;
  assign n257 = x61 ^ x29;
  assign n258 = x61 ^ x28;
  assign n259 = n258 ^ x61;
  assign n260 = x61 ^ x60;
  assign n261 = n260 ^ x61;
  assign n262 = n259 & ~n261;
  assign n263 = n262 ^ x61;
  assign n264 = ~n257 & n263;
  assign n265 = n264 ^ x29;
  assign n266 = n265 ^ x63;
  assign n267 = n266 ^ x63;
  assign n268 = n68 ^ x63;
  assign n269 = n268 ^ x63;
  assign n270 = n267 & ~n269;
  assign n271 = n270 ^ x63;
  assign n274 = n271 ^ x63;
  assign n272 = n271 ^ x62;
  assign n273 = n272 ^ n271;
  assign n275 = n274 ^ n273;
  assign n276 = n271 ^ x30;
  assign n277 = n276 ^ n271;
  assign n278 = n277 ^ n273;
  assign n279 = ~n273 & ~n278;
  assign n280 = n279 ^ n273;
  assign n281 = n275 & ~n280;
  assign n282 = n281 ^ n279;
  assign n283 = n282 ^ n271;
  assign n284 = n283 ^ n273;
  assign n285 = ~n256 & ~n284;
  assign n286 = n285 ^ x31;
  assign n287 = ~n255 & ~n286;
  assign n288 = n159 & n287;
  assign y0 = n288;
endmodule