module Xor(
    input logic a, b//,
    //output logic out
);

    logic c;
    logic d;

    assign c = 0;
    assign d = a;

    //assign out = a ^ b;
    
endmodule
