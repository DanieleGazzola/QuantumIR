module FullAdder(input logic a, b,
                 output logic sum);

    assign sum = a ^ b;
    
endmodule