module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141;
  wire n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272;
  assign n148 = ~x8 & ~x10;
  assign n149 = ~x14 & ~x21;
  assign n150 = n148 & n149;
  assign n151 = ~x13 & n150;
  assign n152 = ~x4 & ~x9;
  assign n153 = ~x12 & n152;
  assign n154 = ~x7 & n153;
  assign n155 = n151 & n154;
  assign n156 = ~x12 & ~x13;
  assign n157 = n156 ^ x9;
  assign n161 = x7 ^ x6;
  assign n158 = ~x6 & ~x7;
  assign n159 = x12 & x13;
  assign n160 = n158 & ~n159;
  assign n162 = n161 ^ n160;
  assign n163 = n162 ^ n160;
  assign n164 = n160 ^ n156;
  assign n165 = n164 ^ n160;
  assign n166 = n163 & n165;
  assign n167 = n166 ^ n160;
  assign n168 = n157 & n167;
  assign n169 = n168 ^ n160;
  assign n170 = n155 & ~n169;
  assign n171 = ~x5 & ~x22;
  assign n172 = ~x11 & n171;
  assign n173 = ~x18 & ~x19;
  assign n174 = ~x16 & n173;
  assign n175 = n172 & n174;
  assign n176 = n170 & n175;
  assign n177 = ~x17 & n176;
  assign n178 = x54 & ~n177;
  assign n179 = ~x0 & ~n178;
  assign n180 = x7 & ~n151;
  assign n182 = x21 ^ x14;
  assign n183 = x14 ^ x13;
  assign n184 = n182 & n183;
  assign n185 = n184 ^ x14;
  assign n186 = n148 & ~n185;
  assign n181 = x10 ^ x8;
  assign n187 = n186 ^ n181;
  assign n188 = n181 ^ x7;
  assign n189 = ~x13 & n149;
  assign n190 = n189 ^ n181;
  assign n191 = ~n181 & ~n190;
  assign n192 = n191 ^ n181;
  assign n193 = ~n188 & ~n192;
  assign n194 = n193 ^ n191;
  assign n195 = n194 ^ n181;
  assign n196 = n195 ^ n189;
  assign n197 = n187 & ~n196;
  assign n198 = n197 ^ n186;
  assign n199 = ~n180 & n198;
  assign n200 = ~x6 & n174;
  assign n201 = n153 & n200;
  assign n202 = n199 & n201;
  assign n203 = ~x17 & x54;
  assign n204 = n172 & n203;
  assign n205 = n202 & n204;
  assign n206 = ~x9 & ~x11;
  assign n207 = n206 ^ n171;
  assign n208 = x54 & ~x56;
  assign n209 = n207 & n208;
  assign n210 = ~n205 & ~n209;
  assign n211 = ~n179 & n210;
  assign n212 = ~x3 & ~x129;
  assign n213 = ~n211 & n212;
  assign n214 = ~n176 & n203;
  assign n215 = ~x1 & n212;
  assign n216 = ~n214 & n215;
  assign n217 = ~x5 & ~n169;
  assign n218 = n203 & n212;
  assign n219 = n174 & n218;
  assign n220 = ~x11 & ~x22;
  assign n221 = ~x4 & n220;
  assign n222 = n150 & n221;
  assign n223 = n219 & n222;
  assign n224 = ~n217 & n223;
  assign n225 = x5 & ~n170;
  assign n226 = n224 & ~n225;
  assign n227 = ~n216 & ~n226;
  assign n228 = ~x42 & ~x44;
  assign n229 = ~x40 & n228;
  assign n230 = ~x38 & ~x50;
  assign n231 = n229 & n230;
  assign n232 = ~x41 & ~x46;
  assign n233 = ~x47 & ~x48;
  assign n234 = n232 & n233;
  assign n235 = ~x43 & n234;
  assign n236 = n231 & n235;
  assign n237 = ~x24 & ~x49;
  assign n238 = ~x45 & n237;
  assign n239 = n236 & n238;
  assign n240 = x82 & ~n239;
  assign n241 = x122 & x127;
  assign n242 = ~x82 & n241;
  assign n243 = ~n240 & ~n242;
  assign n244 = ~x15 & ~x20;
  assign n245 = x82 & ~n244;
  assign n246 = n243 & ~n245;
  assign n247 = x2 & ~n246;
  assign n248 = ~x2 & n244;
  assign n249 = n238 & n248;
  assign n250 = n235 & n249;
  assign n251 = x82 & ~n250;
  assign n252 = x82 & ~n230;
  assign n253 = ~n251 & ~n252;
  assign n254 = x82 & ~n229;
  assign n255 = n253 & ~n254;
  assign n256 = ~n241 & n255;
  assign n257 = ~x65 & n256;
  assign n258 = ~n247 & ~n257;
  assign n259 = ~x129 & ~n258;
  assign n260 = ~x61 & ~x118;
  assign n261 = ~x129 & n260;
  assign n262 = ~n177 & n261;
  assign n263 = ~x123 & ~x129;
  assign n264 = x0 & ~x113;
  assign n265 = n263 & n264;
  assign n266 = ~n262 & ~n265;
  assign n267 = n172 & n218;
  assign n268 = n202 & n267;
  assign n269 = x10 & n268;
  assign n270 = ~x54 & n212;
  assign n271 = x4 & n270;
  assign n272 = ~n269 & ~n271;
  assign n273 = ~x16 & n267;
  assign n274 = n170 & n273;
  assign n275 = ~x29 & ~x59;
  assign n276 = n173 & n275;
  assign n277 = n274 & n276;
  assign n278 = ~x25 & x28;
  assign n279 = n277 & n278;
  assign n280 = x5 & n270;
  assign n281 = ~n279 & ~n280;
  assign n282 = x25 & ~x28;
  assign n283 = n277 & n282;
  assign n284 = x6 & n270;
  assign n285 = ~n283 & ~n284;
  assign n286 = x8 & n268;
  assign n287 = x7 & n270;
  assign n288 = ~n286 & ~n287;
  assign n289 = x21 & n268;
  assign n290 = x8 & n270;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~x5 & n219;
  assign n293 = n170 & n292;
  assign n294 = x11 & ~x22;
  assign n295 = n293 & n294;
  assign n296 = x9 & n270;
  assign n297 = ~n295 & ~n296;
  assign n298 = x14 & n268;
  assign n299 = x10 & n270;
  assign n300 = ~n298 & ~n299;
  assign n301 = n293 ^ n270;
  assign n302 = n301 ^ n270;
  assign n303 = n270 ^ x22;
  assign n304 = n303 ^ n270;
  assign n305 = n302 & n304;
  assign n306 = n305 ^ n270;
  assign n307 = ~x11 & n306;
  assign n308 = n307 ^ n270;
  assign n309 = x18 & ~x19;
  assign n310 = n274 & n309;
  assign n311 = x12 & n270;
  assign n312 = ~n310 & ~n311;
  assign n313 = x29 & x54;
  assign n314 = ~x59 & n313;
  assign n315 = ~x25 & ~x28;
  assign n316 = n314 & n315;
  assign n317 = n212 & n316;
  assign n318 = n177 & n317;
  assign n319 = x13 & n270;
  assign n320 = ~n318 & ~n319;
  assign n321 = x13 & n268;
  assign n322 = x14 & n270;
  assign n323 = ~n321 & ~n322;
  assign n324 = x15 & ~n243;
  assign n326 = ~x70 & ~n241;
  assign n325 = ~x15 & n239;
  assign n327 = n326 ^ n325;
  assign n328 = ~x82 & n327;
  assign n329 = n328 ^ n325;
  assign n330 = ~n324 & ~n329;
  assign n331 = n248 & ~n326;
  assign n332 = ~x129 & ~n331;
  assign n333 = ~n330 & n332;
  assign n334 = x6 & n226;
  assign n335 = x16 & n270;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~x29 & x59;
  assign n338 = n315 & n337;
  assign n339 = n218 & n338;
  assign n340 = n176 & n339;
  assign n341 = x17 & n270;
  assign n342 = ~n340 & ~n341;
  assign n343 = x16 & n173;
  assign n344 = n267 & n343;
  assign n345 = n170 & n344;
  assign n346 = x18 & n270;
  assign n347 = ~n345 & ~n346;
  assign n348 = x54 & n212;
  assign n349 = x17 & n348;
  assign n350 = n176 & n349;
  assign n351 = x19 & n270;
  assign n352 = ~n350 & ~n351;
  assign n353 = n325 ^ x20;
  assign n354 = x82 & ~n353;
  assign n355 = x71 ^ x20;
  assign n356 = n355 ^ x71;
  assign n357 = n356 ^ x82;
  assign n358 = n357 ^ n356;
  assign n361 = ~n241 & ~n355;
  assign n363 = n361 ^ n358;
  assign n359 = n356 ^ x2;
  assign n360 = ~n356 & n359;
  assign n364 = n360 ^ n356;
  assign n365 = ~n363 & ~n364;
  assign n362 = n361 ^ n360;
  assign n366 = n365 ^ n362;
  assign n367 = ~n358 & n366;
  assign n368 = n367 ^ n360;
  assign n369 = n368 ^ n365;
  assign n370 = n369 ^ x20;
  assign n371 = ~x129 & n370;
  assign n372 = ~n354 & n371;
  assign n373 = ~x18 & x19;
  assign n374 = n274 & n373;
  assign n375 = x21 & n270;
  assign n376 = ~n374 & ~n375;
  assign n377 = n170 & n224;
  assign n378 = x22 & n270;
  assign n379 = ~n377 & ~n378;
  assign n380 = ~x23 & x55;
  assign n381 = x61 & ~x129;
  assign n382 = ~n380 & n381;
  assign n383 = x63 & n256;
  assign n386 = x82 & ~n249;
  assign n387 = n241 & ~n386;
  assign n384 = x82 & n236;
  assign n385 = ~x45 & n384;
  assign n388 = n387 ^ n385;
  assign n389 = n388 ^ n385;
  assign n390 = x82 & ~n385;
  assign n391 = n390 ^ n385;
  assign n392 = n391 ^ n385;
  assign n393 = ~n389 & ~n392;
  assign n394 = n393 ^ n385;
  assign n395 = ~x24 & ~n394;
  assign n396 = n395 ^ n385;
  assign n397 = ~x129 & ~n396;
  assign n398 = ~n383 & n397;
  assign n399 = ~x26 & ~x27;
  assign n404 = x53 & x58;
  assign n405 = ~x85 & ~n404;
  assign n400 = ~x53 & ~x58;
  assign n406 = n405 ^ n400;
  assign n401 = ~x85 & n400;
  assign n402 = x26 & x27;
  assign n403 = n401 & ~n402;
  assign n407 = n406 ^ n403;
  assign n408 = n399 & n407;
  assign n409 = n408 ^ n403;
  assign n410 = ~x116 & n409;
  assign n411 = ~x95 & ~x100;
  assign n412 = ~x97 & n411;
  assign n413 = ~x110 & ~n412;
  assign n414 = n399 & n401;
  assign n415 = n413 & n414;
  assign n416 = ~x39 & ~x52;
  assign n417 = ~x51 & n416;
  assign n418 = x26 & x116;
  assign n419 = n417 & n418;
  assign n420 = n403 & ~n419;
  assign n421 = ~n415 & n420;
  assign n422 = ~n410 & ~n421;
  assign n423 = x27 & x116;
  assign n424 = ~n417 & n423;
  assign n425 = n212 & ~n424;
  assign n426 = x116 & ~n399;
  assign n427 = ~x25 & ~n426;
  assign n428 = n425 & ~n427;
  assign n429 = ~n422 & n428;
  assign n430 = ~x96 & ~x110;
  assign n431 = n430 ^ x116;
  assign n432 = ~x85 & n431;
  assign n433 = n432 ^ x116;
  assign n434 = x100 & n433;
  assign n435 = n212 & n399;
  assign n436 = n400 & n435;
  assign n437 = n434 & n436;
  assign n438 = ~n429 & ~n437;
  assign n439 = x116 & n417;
  assign n440 = n401 & ~n439;
  assign n441 = x26 & ~x27;
  assign n442 = n212 & n441;
  assign n443 = n440 & n442;
  assign n444 = ~n437 & ~n443;
  assign n445 = ~x26 & x27;
  assign n446 = n440 & n445;
  assign n447 = x85 & x116;
  assign n448 = ~x95 & ~n447;
  assign n449 = n399 & n400;
  assign n450 = ~n448 & n449;
  assign n451 = ~x100 & n450;
  assign n452 = n433 & n451;
  assign n453 = ~n446 & ~n452;
  assign n454 = n212 & ~n453;
  assign n455 = ~x26 & x28;
  assign n456 = ~n413 & n455;
  assign n457 = ~n419 & ~n456;
  assign n458 = ~x27 & n401;
  assign n459 = ~n457 & n458;
  assign n460 = n454 ^ n410;
  assign n461 = n460 ^ n454;
  assign n462 = n454 ^ x28;
  assign n463 = n461 & n462;
  assign n464 = n463 ^ n454;
  assign n465 = ~n459 & ~n464;
  assign n466 = n212 & ~n465;
  assign n467 = ~n413 & n414;
  assign n468 = ~n410 & ~n467;
  assign n469 = x29 & ~n468;
  assign n470 = x53 & x116;
  assign n471 = n405 & ~n470;
  assign n472 = n435 & n471;
  assign n473 = ~x53 & x97;
  assign n474 = n411 & n430;
  assign n475 = n474 ^ x116;
  assign n476 = x116 ^ x58;
  assign n477 = n476 ^ x116;
  assign n478 = n477 ^ n473;
  assign n479 = n475 & ~n478;
  assign n480 = n479 ^ n474;
  assign n481 = n473 & n480;
  assign n482 = n481 ^ x53;
  assign n483 = n472 & n482;
  assign n484 = ~n410 & n483;
  assign n485 = ~n469 & ~n484;
  assign n486 = n212 & ~n485;
  assign n487 = x106 ^ x88;
  assign n488 = n487 ^ x88;
  assign n489 = x60 ^ x30;
  assign n490 = x109 & n489;
  assign n491 = n490 ^ x30;
  assign n492 = n491 ^ x88;
  assign n493 = ~n488 & n492;
  assign n494 = n493 ^ x88;
  assign n495 = ~x129 & n494;
  assign n496 = x106 ^ x89;
  assign n497 = n496 ^ x89;
  assign n498 = x31 ^ x30;
  assign n499 = ~x109 & n498;
  assign n500 = n499 ^ x30;
  assign n501 = n500 ^ x89;
  assign n502 = ~n497 & n501;
  assign n503 = n502 ^ x89;
  assign n504 = ~x129 & n503;
  assign n505 = x106 ^ x99;
  assign n506 = n505 ^ x99;
  assign n507 = x32 ^ x31;
  assign n508 = ~x109 & n507;
  assign n509 = n508 ^ x31;
  assign n510 = n509 ^ x99;
  assign n511 = ~n506 & n510;
  assign n512 = n511 ^ x99;
  assign n513 = ~x129 & n512;
  assign n514 = x106 ^ x90;
  assign n515 = n514 ^ x90;
  assign n516 = x33 ^ x32;
  assign n517 = ~x109 & n516;
  assign n518 = n517 ^ x32;
  assign n519 = n518 ^ x90;
  assign n520 = ~n515 & n519;
  assign n521 = n520 ^ x90;
  assign n522 = ~x129 & n521;
  assign n523 = x106 ^ x91;
  assign n524 = n523 ^ x91;
  assign n525 = x34 ^ x33;
  assign n526 = ~x109 & n525;
  assign n527 = n526 ^ x33;
  assign n528 = n527 ^ x91;
  assign n529 = ~n524 & n528;
  assign n530 = n529 ^ x91;
  assign n531 = ~x129 & n530;
  assign n532 = x106 ^ x92;
  assign n533 = n532 ^ x92;
  assign n534 = x35 ^ x34;
  assign n535 = ~x109 & n534;
  assign n536 = n535 ^ x34;
  assign n537 = n536 ^ x92;
  assign n538 = ~n533 & n537;
  assign n539 = n538 ^ x92;
  assign n540 = ~x129 & n539;
  assign n541 = x106 ^ x98;
  assign n542 = n541 ^ x98;
  assign n543 = x36 ^ x35;
  assign n544 = ~x109 & n543;
  assign n545 = n544 ^ x35;
  assign n546 = n545 ^ x98;
  assign n547 = ~n542 & n546;
  assign n548 = n547 ^ x98;
  assign n549 = ~x129 & n548;
  assign n550 = x106 ^ x93;
  assign n551 = n550 ^ x93;
  assign n552 = x37 ^ x36;
  assign n553 = ~x109 & n552;
  assign n554 = n553 ^ x36;
  assign n555 = n554 ^ x93;
  assign n556 = ~n551 & n555;
  assign n557 = n556 ^ x93;
  assign n558 = ~x129 & n557;
  assign n559 = x74 ^ x38;
  assign n560 = ~n241 & ~n559;
  assign n561 = n560 ^ x38;
  assign n562 = n253 & ~n561;
  assign n563 = n229 ^ x38;
  assign n564 = x82 & ~n563;
  assign n565 = ~x129 & ~n564;
  assign n566 = ~n562 & n565;
  assign n567 = ~x51 & x109;
  assign n568 = ~x52 & n567;
  assign n569 = n568 ^ x39;
  assign n570 = ~x106 & ~n569;
  assign n571 = ~x129 & ~n570;
  assign n572 = ~x73 & ~n241;
  assign n573 = n253 & ~n572;
  assign n574 = ~n254 & ~n573;
  assign n575 = x82 & ~n228;
  assign n576 = ~n242 & ~n575;
  assign n577 = x40 & ~n576;
  assign n578 = ~n574 & ~n577;
  assign n579 = ~x129 & ~n578;
  assign n580 = ~x46 & n231;
  assign n581 = n580 ^ x41;
  assign n582 = x82 & ~n581;
  assign n583 = ~x129 & ~n582;
  assign n584 = x76 ^ x41;
  assign n585 = ~n241 & ~n584;
  assign n586 = n585 ^ x41;
  assign n587 = ~n251 & ~n586;
  assign n588 = n583 & ~n587;
  assign n589 = n228 & ~n255;
  assign n590 = x44 & x82;
  assign n591 = ~n242 & ~n590;
  assign n592 = x42 & ~n591;
  assign n593 = ~x72 & ~n241;
  assign n594 = ~n575 & n593;
  assign n595 = ~n592 & ~n594;
  assign n596 = ~n589 & n595;
  assign n597 = ~x129 & ~n596;
  assign n598 = n231 & n232;
  assign n599 = n598 ^ x43;
  assign n600 = x82 & ~n599;
  assign n601 = ~x129 & ~n600;
  assign n602 = x77 ^ x43;
  assign n603 = ~n241 & ~n602;
  assign n604 = n603 ^ x43;
  assign n605 = ~n251 & ~n604;
  assign n606 = n601 & ~n605;
  assign n607 = x67 ^ x44;
  assign n608 = ~n241 & ~n607;
  assign n609 = n608 ^ x44;
  assign n610 = n255 & ~n609;
  assign n611 = ~x129 & ~n590;
  assign n612 = ~n610 & n611;
  assign n613 = ~x68 & ~n241;
  assign n614 = ~n386 & ~n613;
  assign n615 = ~n390 & ~n614;
  assign n616 = ~x82 & ~n241;
  assign n617 = x45 & ~n616;
  assign n618 = ~n384 & n617;
  assign n619 = ~n615 & ~n618;
  assign n620 = ~x129 & ~n619;
  assign n621 = x75 ^ x46;
  assign n622 = ~n241 & ~n621;
  assign n623 = n622 ^ x46;
  assign n624 = n255 & ~n623;
  assign n625 = n231 ^ x46;
  assign n626 = x82 & ~n625;
  assign n627 = ~x129 & ~n626;
  assign n628 = ~n624 & n627;
  assign n629 = ~x43 & n598;
  assign n630 = n629 ^ x47;
  assign n631 = x82 & ~n630;
  assign n632 = x64 ^ x47;
  assign n633 = ~n241 & ~n632;
  assign n634 = n633 ^ x47;
  assign n635 = ~n251 & ~n634;
  assign n636 = ~x129 & ~n635;
  assign n637 = ~n631 & n636;
  assign n638 = ~x47 & n629;
  assign n639 = n638 ^ x48;
  assign n640 = x82 & ~n639;
  assign n641 = x48 & ~n616;
  assign n642 = ~x62 & ~n241;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n386 & n643;
  assign n645 = ~x129 & ~n644;
  assign n646 = ~n640 & n645;
  assign n647 = ~x24 & n385;
  assign n648 = x49 & ~n616;
  assign n649 = ~n647 & n648;
  assign n650 = x82 & ~n248;
  assign n651 = ~x69 & ~n241;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n240 & ~n652;
  assign n654 = ~n649 & ~n653;
  assign n655 = ~x129 & ~n654;
  assign n656 = ~x66 & ~n241;
  assign n657 = n250 & ~n656;
  assign n658 = ~n242 & ~n252;
  assign n659 = ~n254 & n658;
  assign n660 = ~n657 & n659;
  assign n661 = ~x50 & ~n660;
  assign n662 = ~x38 & n229;
  assign n663 = n252 & n662;
  assign n664 = x66 & n616;
  assign n665 = ~x129 & ~n664;
  assign n666 = ~n663 & n665;
  assign n667 = ~n661 & n666;
  assign n668 = x109 ^ x51;
  assign n669 = ~x106 & ~n668;
  assign n670 = ~x129 & ~n669;
  assign n671 = n567 ^ x52;
  assign n672 = ~x106 & ~n671;
  assign n673 = ~x129 & ~n672;
  assign n674 = ~x129 & ~n256;
  assign n675 = x114 & ~x122;
  assign n676 = n263 & n675;
  assign n677 = n399 & n406;
  assign n678 = ~n403 & ~n677;
  assign n679 = n212 & ~n678;
  assign n680 = ~x37 & ~x58;
  assign n681 = n680 ^ x94;
  assign n682 = x58 & ~x116;
  assign n683 = n682 ^ n680;
  assign n684 = n680 ^ n418;
  assign n685 = ~n680 & n684;
  assign n686 = n685 ^ n680;
  assign n687 = ~n683 & ~n686;
  assign n688 = n687 ^ n685;
  assign n689 = n688 ^ n680;
  assign n690 = n689 ^ n418;
  assign n691 = ~n681 & n690;
  assign n692 = n691 ^ x94;
  assign n693 = n679 & n692;
  assign n694 = x58 & x116;
  assign n695 = x60 ^ x57;
  assign n696 = n694 & n695;
  assign n697 = n696 ^ x57;
  assign n698 = n679 & n697;
  assign n699 = n417 & n426;
  assign n700 = ~n682 & ~n699;
  assign n701 = n679 & ~n700;
  assign n702 = x59 & ~n468;
  assign n703 = x96 & n415;
  assign n704 = ~n702 & ~n703;
  assign n705 = n212 & ~n704;
  assign n706 = ~x117 & ~x122;
  assign n707 = x123 ^ x60;
  assign n708 = n706 & n707;
  assign n709 = n708 ^ x60;
  assign n710 = ~x114 & ~x122;
  assign n711 = x123 & ~x129;
  assign n712 = n710 & n711;
  assign n713 = x132 & x133;
  assign n714 = x131 & n713;
  assign n715 = ~x138 & n714;
  assign n716 = x136 & ~x137;
  assign n717 = n715 & n716;
  assign n718 = n717 ^ x62;
  assign n719 = n718 ^ x62;
  assign n720 = x140 ^ x62;
  assign n721 = n719 & ~n720;
  assign n722 = n721 ^ x62;
  assign n723 = ~x129 & n722;
  assign n724 = n717 ^ x63;
  assign n725 = n724 ^ x63;
  assign n726 = x142 ^ x63;
  assign n727 = n725 & ~n726;
  assign n728 = n727 ^ x63;
  assign n729 = ~x129 & n728;
  assign n730 = n717 ^ x64;
  assign n731 = n730 ^ x64;
  assign n732 = x139 ^ x64;
  assign n733 = n731 & ~n732;
  assign n734 = n733 ^ x64;
  assign n735 = ~x129 & n734;
  assign n736 = n717 ^ x65;
  assign n737 = n736 ^ x65;
  assign n738 = x146 ^ x65;
  assign n739 = n737 & ~n738;
  assign n740 = n739 ^ x65;
  assign n741 = ~x129 & n740;
  assign n742 = ~x136 & ~x137;
  assign n743 = n715 & n742;
  assign n744 = n743 ^ x66;
  assign n745 = n744 ^ x66;
  assign n746 = x143 ^ x66;
  assign n747 = n745 & ~n746;
  assign n748 = n747 ^ x66;
  assign n749 = ~x129 & n748;
  assign n750 = n743 ^ x67;
  assign n751 = n750 ^ x67;
  assign n752 = x139 ^ x67;
  assign n753 = n751 & ~n752;
  assign n754 = n753 ^ x67;
  assign n755 = ~x129 & n754;
  assign n756 = n717 ^ x68;
  assign n757 = n756 ^ x68;
  assign n758 = x141 ^ x68;
  assign n759 = n757 & ~n758;
  assign n760 = n759 ^ x68;
  assign n761 = ~x129 & n760;
  assign n762 = n717 ^ x69;
  assign n763 = n762 ^ x69;
  assign n764 = x143 ^ x69;
  assign n765 = n763 & ~n764;
  assign n766 = n765 ^ x69;
  assign n767 = ~x129 & n766;
  assign n768 = n717 ^ x70;
  assign n769 = n768 ^ x70;
  assign n770 = x144 ^ x70;
  assign n771 = n769 & ~n770;
  assign n772 = n771 ^ x70;
  assign n773 = ~x129 & n772;
  assign n774 = n717 ^ x71;
  assign n775 = n774 ^ x71;
  assign n776 = x145 ^ x71;
  assign n777 = n775 & ~n776;
  assign n778 = n777 ^ x71;
  assign n779 = ~x129 & n778;
  assign n780 = n743 ^ x72;
  assign n781 = n780 ^ x72;
  assign n782 = x140 ^ x72;
  assign n783 = n781 & ~n782;
  assign n784 = n783 ^ x72;
  assign n785 = ~x129 & n784;
  assign n786 = n743 ^ x73;
  assign n787 = n786 ^ x73;
  assign n788 = x141 ^ x73;
  assign n789 = n787 & ~n788;
  assign n790 = n789 ^ x73;
  assign n791 = ~x129 & n790;
  assign n792 = n743 ^ x74;
  assign n793 = n792 ^ x74;
  assign n794 = x142 ^ x74;
  assign n795 = n793 & ~n794;
  assign n796 = n795 ^ x74;
  assign n797 = ~x129 & n796;
  assign n798 = n743 ^ x75;
  assign n799 = n798 ^ x75;
  assign n800 = x144 ^ x75;
  assign n801 = n799 & ~n800;
  assign n802 = n801 ^ x75;
  assign n803 = ~x129 & n802;
  assign n804 = n743 ^ x76;
  assign n805 = n804 ^ x76;
  assign n806 = x145 ^ x76;
  assign n807 = n805 & ~n806;
  assign n808 = n807 ^ x76;
  assign n809 = ~x129 & n808;
  assign n810 = n743 ^ x77;
  assign n811 = n810 ^ x77;
  assign n812 = x146 ^ x77;
  assign n813 = n811 & ~n812;
  assign n814 = n813 ^ x77;
  assign n815 = ~x129 & n814;
  assign n816 = ~x136 & x137;
  assign n817 = n715 & n816;
  assign n818 = n817 ^ x78;
  assign n819 = n818 ^ x78;
  assign n820 = x142 ^ x78;
  assign n821 = n819 & n820;
  assign n822 = n821 ^ x78;
  assign n823 = ~x129 & n822;
  assign n824 = n817 ^ x79;
  assign n825 = n824 ^ x79;
  assign n826 = x143 ^ x79;
  assign n827 = n825 & n826;
  assign n828 = n827 ^ x79;
  assign n829 = ~x129 & n828;
  assign n830 = n817 ^ x80;
  assign n831 = n830 ^ x80;
  assign n832 = x144 ^ x80;
  assign n833 = n831 & n832;
  assign n834 = n833 ^ x80;
  assign n835 = ~x129 & n834;
  assign n836 = n817 ^ x81;
  assign n837 = n836 ^ x81;
  assign n838 = x145 ^ x81;
  assign n839 = n837 & n838;
  assign n840 = n839 ^ x81;
  assign n841 = ~x129 & n840;
  assign n842 = n817 ^ x82;
  assign n843 = n842 ^ x82;
  assign n844 = x146 ^ x82;
  assign n845 = n843 & n844;
  assign n846 = n845 ^ x82;
  assign n847 = ~x129 & n846;
  assign n861 = x138 ^ x115;
  assign n862 = n861 ^ x115;
  assign n863 = x115 ^ x87;
  assign n864 = ~n862 & ~n863;
  assign n865 = n864 ^ x115;
  assign n866 = n865 ^ x137;
  assign n867 = n866 ^ n865;
  assign n868 = x138 ^ x119;
  assign n869 = n868 ^ x119;
  assign n870 = x119 ^ x72;
  assign n871 = ~n869 & ~n870;
  assign n872 = n871 ^ x119;
  assign n873 = n872 ^ n865;
  assign n874 = ~n867 & ~n873;
  assign n875 = n874 ^ n865;
  assign n848 = x62 ^ x31;
  assign n849 = ~x137 & ~n848;
  assign n850 = n849 ^ x31;
  assign n851 = n850 ^ x138;
  assign n852 = n851 ^ n850;
  assign n853 = n852 ^ x136;
  assign n854 = x137 ^ x89;
  assign n855 = ~x137 & ~n854;
  assign n856 = n855 ^ n850;
  assign n857 = n856 ^ x137;
  assign n858 = n853 & ~n857;
  assign n859 = n858 ^ n855;
  assign n860 = n859 ^ x137;
  assign n876 = n875 ^ n860;
  assign n877 = ~x136 & n876;
  assign n878 = n877 ^ n860;
  assign n879 = n817 ^ x84;
  assign n880 = n879 ^ x84;
  assign n881 = x141 ^ x84;
  assign n882 = n880 & n881;
  assign n883 = n882 ^ x84;
  assign n884 = ~x129 & n883;
  assign n885 = x116 ^ x85;
  assign n886 = n885 ^ x116;
  assign n887 = x96 & n413;
  assign n888 = n887 ^ x116;
  assign n889 = ~n886 & ~n888;
  assign n890 = n889 ^ x116;
  assign n891 = n436 & ~n890;
  assign n892 = n817 ^ x86;
  assign n893 = n892 ^ x86;
  assign n894 = x139 ^ x86;
  assign n895 = n893 & n894;
  assign n896 = n895 ^ x86;
  assign n897 = ~x129 & n896;
  assign n898 = n817 ^ x87;
  assign n899 = n898 ^ x87;
  assign n900 = x140 ^ x87;
  assign n901 = n899 & n900;
  assign n902 = n901 ^ x87;
  assign n903 = ~x129 & n902;
  assign n904 = x136 & x137;
  assign n905 = n715 & n904;
  assign n906 = n905 ^ x88;
  assign n907 = n906 ^ x88;
  assign n908 = x139 ^ x88;
  assign n909 = n907 & n908;
  assign n910 = n909 ^ x88;
  assign n911 = ~x129 & n910;
  assign n912 = n905 ^ x89;
  assign n913 = n912 ^ x89;
  assign n914 = x140 ^ x89;
  assign n915 = n913 & n914;
  assign n916 = n915 ^ x89;
  assign n917 = ~x129 & n916;
  assign n918 = n905 ^ x90;
  assign n919 = n918 ^ x90;
  assign n920 = x142 ^ x90;
  assign n921 = n919 & n920;
  assign n922 = n921 ^ x90;
  assign n923 = ~x129 & n922;
  assign n924 = n905 ^ x91;
  assign n925 = n924 ^ x91;
  assign n926 = x143 ^ x91;
  assign n927 = n925 & n926;
  assign n928 = n927 ^ x91;
  assign n929 = ~x129 & n928;
  assign n930 = n905 ^ x92;
  assign n931 = n930 ^ x92;
  assign n932 = x144 ^ x92;
  assign n933 = n931 & n932;
  assign n934 = n933 ^ x92;
  assign n935 = ~x129 & n934;
  assign n936 = n905 ^ x93;
  assign n937 = n936 ^ x93;
  assign n938 = x146 ^ x93;
  assign n939 = n937 & n938;
  assign n940 = n939 ^ x93;
  assign n941 = ~x129 & n940;
  assign n942 = x82 & x138;
  assign n943 = n742 & n942;
  assign n944 = n714 & n943;
  assign n945 = n944 ^ x94;
  assign n946 = n945 ^ x94;
  assign n947 = x142 ^ x94;
  assign n948 = n946 & n947;
  assign n949 = n948 ^ x94;
  assign n950 = ~x129 & n949;
  assign n951 = ~x3 & ~x110;
  assign n952 = ~n714 & ~n951;
  assign n953 = n952 ^ x143;
  assign n954 = n953 ^ x143;
  assign n955 = x143 ^ x95;
  assign n956 = n955 ^ x143;
  assign n957 = ~n954 & n956;
  assign n958 = n957 ^ x143;
  assign n959 = ~n944 & n958;
  assign n960 = n959 ^ x143;
  assign n961 = ~x129 & n960;
  assign n962 = n952 ^ x146;
  assign n963 = n962 ^ x146;
  assign n964 = x146 ^ x96;
  assign n965 = n964 ^ x146;
  assign n966 = ~n963 & n965;
  assign n967 = n966 ^ x146;
  assign n968 = ~n944 & n967;
  assign n969 = n968 ^ x146;
  assign n970 = ~x129 & n969;
  assign n971 = n952 ^ x145;
  assign n972 = n971 ^ x145;
  assign n973 = x145 ^ x97;
  assign n974 = n973 ^ x145;
  assign n975 = ~n972 & n974;
  assign n976 = n975 ^ x145;
  assign n977 = ~n944 & n976;
  assign n978 = n977 ^ x145;
  assign n979 = ~x129 & n978;
  assign n980 = n905 ^ x98;
  assign n981 = n980 ^ x98;
  assign n982 = x145 ^ x98;
  assign n983 = n981 & n982;
  assign n984 = n983 ^ x98;
  assign n985 = ~x129 & n984;
  assign n986 = n905 ^ x99;
  assign n987 = n986 ^ x99;
  assign n988 = x141 ^ x99;
  assign n989 = n987 & n988;
  assign n990 = n989 ^ x99;
  assign n991 = ~x129 & n990;
  assign n992 = n952 ^ x144;
  assign n993 = n992 ^ x144;
  assign n994 = x144 ^ x100;
  assign n995 = n994 ^ x144;
  assign n996 = ~n993 & n995;
  assign n997 = n996 ^ x144;
  assign n998 = ~n944 & n997;
  assign n999 = n998 ^ x144;
  assign n1000 = ~x129 & n999;
  assign n1001 = ~x65 & n716;
  assign n1002 = ~x138 & ~n1001;
  assign n1003 = x136 ^ x82;
  assign n1004 = n1003 ^ x82;
  assign n1005 = x82 ^ x37;
  assign n1006 = n1004 & n1005;
  assign n1007 = n1006 ^ x82;
  assign n1008 = x137 & n1007;
  assign n1009 = n1002 & ~n1008;
  assign n1010 = x137 ^ x136;
  assign n1011 = n1010 ^ x138;
  assign n1012 = x137 ^ x96;
  assign n1013 = n1012 ^ x96;
  assign n1014 = x96 ^ x93;
  assign n1015 = ~n1013 & n1014;
  assign n1016 = n1015 ^ x96;
  assign n1017 = n1016 ^ n1010;
  assign n1018 = n1011 & n1017;
  assign n1019 = n1018 ^ n1015;
  assign n1020 = n1019 ^ x96;
  assign n1021 = n1020 ^ x138;
  assign n1022 = n1010 & n1021;
  assign n1023 = n1022 ^ n1010;
  assign n1024 = n1023 ^ x138;
  assign n1025 = ~n1009 & ~n1024;
  assign n1026 = x138 ^ x124;
  assign n1027 = n1026 ^ x124;
  assign n1028 = x124 ^ x77;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = n1029 ^ x124;
  assign n1031 = n742 & n1030;
  assign n1032 = ~n1025 & ~n1031;
  assign n1033 = x136 ^ x69;
  assign n1034 = n1033 ^ x69;
  assign n1035 = x69 ^ x66;
  assign n1036 = ~n1034 & n1035;
  assign n1037 = n1036 ^ x69;
  assign n1038 = ~x137 & ~n1037;
  assign n1039 = x138 ^ x137;
  assign n1040 = x136 ^ x34;
  assign n1041 = n1040 ^ x34;
  assign n1042 = x79 ^ x34;
  assign n1043 = ~n1041 & n1042;
  assign n1044 = n1043 ^ x34;
  assign n1045 = n1044 ^ x138;
  assign n1046 = ~n1039 & ~n1045;
  assign n1047 = n1046 ^ n1043;
  assign n1048 = n1047 ^ x34;
  assign n1049 = n1048 ^ x137;
  assign n1050 = ~x138 & n1049;
  assign n1051 = n1050 ^ x138;
  assign n1052 = n1051 ^ x138;
  assign n1053 = ~n1038 & n1052;
  assign n1054 = x137 ^ x95;
  assign n1055 = n1054 ^ x95;
  assign n1056 = x95 ^ x91;
  assign n1057 = ~n1055 & n1056;
  assign n1058 = n1057 ^ x95;
  assign n1059 = n1058 ^ n1010;
  assign n1060 = n1011 & n1059;
  assign n1061 = n1060 ^ n1057;
  assign n1062 = n1061 ^ x95;
  assign n1063 = n1062 ^ x138;
  assign n1064 = n1010 & n1063;
  assign n1065 = n1064 ^ n1010;
  assign n1066 = n1065 ^ x138;
  assign n1067 = ~n1053 & ~n1066;
  assign n1068 = x78 & n816;
  assign n1069 = ~x138 & ~n1068;
  assign n1070 = x137 ^ x63;
  assign n1071 = n1070 ^ x63;
  assign n1072 = x63 ^ x33;
  assign n1073 = n1071 & ~n1072;
  assign n1074 = n1073 ^ x63;
  assign n1075 = n1074 ^ x74;
  assign n1076 = n1075 ^ n1074;
  assign n1077 = n1074 ^ x137;
  assign n1078 = n1077 ^ n1074;
  assign n1079 = ~n1076 & ~n1078;
  assign n1080 = n1079 ^ n1074;
  assign n1081 = ~x136 & ~n1080;
  assign n1082 = n1081 ^ n1074;
  assign n1083 = n1069 & n1082;
  assign n1084 = x137 ^ x94;
  assign n1085 = n1084 ^ x94;
  assign n1086 = x94 ^ x90;
  assign n1087 = ~n1085 & n1086;
  assign n1088 = n1087 ^ x94;
  assign n1089 = n1088 ^ n1010;
  assign n1090 = n1011 & n1089;
  assign n1091 = n1090 ^ n1087;
  assign n1092 = n1091 ^ x94;
  assign n1093 = n1092 ^ x138;
  assign n1094 = n1010 & n1093;
  assign n1095 = n1094 ^ n1010;
  assign n1096 = n1095 ^ x138;
  assign n1097 = ~n1083 & ~n1096;
  assign n1098 = x136 ^ x68;
  assign n1099 = n1098 ^ x68;
  assign n1100 = x73 ^ x68;
  assign n1101 = ~n1099 & n1100;
  assign n1102 = n1101 ^ x68;
  assign n1103 = n1102 ^ x138;
  assign n1104 = n1039 & n1103;
  assign n1105 = n1104 ^ n1101;
  assign n1106 = n1105 ^ x68;
  assign n1107 = n1106 ^ x137;
  assign n1108 = ~x138 & n1107;
  assign n1109 = n1108 ^ x138;
  assign n1110 = n1109 ^ x138;
  assign n1111 = x136 ^ x84;
  assign n1112 = n1111 ^ x84;
  assign n1113 = x84 ^ x32;
  assign n1114 = n1112 & n1113;
  assign n1115 = n1114 ^ x84;
  assign n1116 = x137 & n1115;
  assign n1117 = n1110 & ~n1116;
  assign n1118 = x137 ^ x112;
  assign n1119 = n1118 ^ x112;
  assign n1120 = x112 ^ x99;
  assign n1121 = ~n1119 & ~n1120;
  assign n1122 = n1121 ^ x112;
  assign n1123 = n1122 ^ n1010;
  assign n1124 = n1011 & ~n1123;
  assign n1125 = n1124 ^ n1121;
  assign n1126 = n1125 ^ x112;
  assign n1127 = n1126 ^ x138;
  assign n1128 = n1010 & ~n1127;
  assign n1129 = n1128 ^ n1010;
  assign n1130 = n1129 ^ x138;
  assign n1131 = ~n1117 & ~n1130;
  assign n1145 = x137 ^ x125;
  assign n1146 = n1145 ^ x125;
  assign n1147 = x125 ^ x100;
  assign n1148 = n1146 & n1147;
  assign n1149 = n1148 ^ x125;
  assign n1150 = n1149 ^ x92;
  assign n1151 = n1150 ^ n1149;
  assign n1152 = n1149 ^ x137;
  assign n1153 = n1152 ^ n1149;
  assign n1154 = n1151 & ~n1153;
  assign n1155 = n1154 ^ n1149;
  assign n1156 = x136 & n1155;
  assign n1157 = n1156 ^ n1149;
  assign n1137 = x137 ^ x80;
  assign n1138 = n1137 ^ x80;
  assign n1139 = x80 ^ x75;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = n1140 ^ x80;
  assign n1132 = x137 ^ x70;
  assign n1133 = n1132 ^ x70;
  assign n1134 = x70 ^ x35;
  assign n1135 = n1133 & ~n1134;
  assign n1136 = n1135 ^ x70;
  assign n1142 = n1141 ^ n1136;
  assign n1143 = x136 & ~n1142;
  assign n1144 = n1143 ^ n1141;
  assign n1158 = n1157 ^ n1144;
  assign n1159 = x138 & n1158;
  assign n1160 = n1159 ^ n1144;
  assign n1161 = ~n415 & ~n447;
  assign n1162 = n212 & ~n1161;
  assign n1178 = x71 ^ x36;
  assign n1179 = ~x137 & ~n1178;
  assign n1180 = n1179 ^ x36;
  assign n1181 = n1180 ^ x137;
  assign n1182 = n1181 ^ n1180;
  assign n1183 = n1180 ^ x98;
  assign n1184 = n1183 ^ n1180;
  assign n1185 = ~n1182 & n1184;
  assign n1186 = n1185 ^ n1180;
  assign n1187 = x138 & n1186;
  assign n1188 = n1187 ^ n1180;
  assign n1163 = x138 ^ x76;
  assign n1164 = n1163 ^ x76;
  assign n1165 = x76 ^ x23;
  assign n1166 = n1164 & ~n1165;
  assign n1167 = n1166 ^ x76;
  assign n1168 = n1167 ^ x137;
  assign n1169 = n1168 ^ n1167;
  assign n1170 = x138 ^ x97;
  assign n1171 = n1170 ^ x97;
  assign n1172 = x97 ^ x81;
  assign n1173 = ~n1171 & n1172;
  assign n1174 = n1173 ^ x97;
  assign n1175 = n1174 ^ n1167;
  assign n1176 = n1169 & ~n1175;
  assign n1177 = n1176 ^ n1167;
  assign n1189 = n1188 ^ n1177;
  assign n1190 = ~x136 & ~n1189;
  assign n1191 = n1190 ^ n1188;
  assign n1205 = x138 ^ x120;
  assign n1206 = n1205 ^ x120;
  assign n1207 = x120 ^ x67;
  assign n1208 = ~n1206 & ~n1207;
  assign n1209 = n1208 ^ x120;
  assign n1210 = n1209 ^ x137;
  assign n1211 = n1210 ^ n1209;
  assign n1212 = x138 ^ x111;
  assign n1213 = n1212 ^ x111;
  assign n1214 = x111 ^ x86;
  assign n1215 = ~n1213 & n1214;
  assign n1216 = n1215 ^ x111;
  assign n1217 = n1216 ^ n1209;
  assign n1218 = n1211 & n1217;
  assign n1219 = n1218 ^ n1209;
  assign n1192 = x64 ^ x30;
  assign n1193 = ~x137 & ~n1192;
  assign n1194 = n1193 ^ x30;
  assign n1195 = n1194 ^ x138;
  assign n1196 = n1195 ^ n1194;
  assign n1197 = n1196 ^ x136;
  assign n1198 = x137 ^ x88;
  assign n1199 = ~x137 & ~n1198;
  assign n1200 = n1199 ^ n1194;
  assign n1201 = n1200 ^ x137;
  assign n1202 = n1197 & ~n1201;
  assign n1203 = n1202 ^ n1199;
  assign n1204 = n1203 ^ x137;
  assign n1220 = n1219 ^ n1204;
  assign n1221 = ~x136 & ~n1220;
  assign n1222 = n1221 ^ n1204;
  assign n1223 = ~n417 & n445;
  assign n1224 = ~n441 & ~n1223;
  assign n1225 = x116 & n212;
  assign n1226 = ~n1224 & n1225;
  assign n1227 = x58 ^ x53;
  assign n1228 = ~n473 & n1227;
  assign n1229 = n1225 & n1228;
  assign n1230 = ~x129 & n714;
  assign n1231 = n943 ^ x139;
  assign n1232 = n1231 ^ x139;
  assign n1233 = x139 ^ x111;
  assign n1234 = ~n1232 & n1233;
  assign n1235 = n1234 ^ x139;
  assign n1236 = n1230 & n1235;
  assign n1237 = n943 ^ x141;
  assign n1238 = n1237 ^ x141;
  assign n1239 = x141 ^ x112;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = n1240 ^ x141;
  assign n1242 = n1230 & n1241;
  assign n1243 = x113 ^ x54;
  assign n1244 = n1243 ^ x113;
  assign n1245 = n220 ^ x113;
  assign n1246 = n1244 & n1245;
  assign n1247 = n1246 ^ x113;
  assign n1248 = n212 & ~n1247;
  assign n1249 = n943 ^ x140;
  assign n1250 = n1249 ^ x140;
  assign n1251 = x140 ^ x115;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = n1252 ^ x140;
  assign n1254 = n1230 & n1253;
  assign n1255 = ~n154 & n348;
  assign n1256 = x122 & ~x129;
  assign n1257 = ~x54 & x118;
  assign n1258 = ~n316 & ~n1257;
  assign n1259 = ~x129 & ~n1258;
  assign n1260 = ~x129 & ~n411;
  assign n1261 = ~x120 & n951;
  assign n1262 = ~x111 & ~x129;
  assign n1263 = ~n1261 & n1262;
  assign n1264 = x81 & x120;
  assign n1265 = ~x129 & n1264;
  assign n1266 = ~x129 & ~x134;
  assign n1267 = ~x129 & ~x135;
  assign n1268 = x57 & ~x129;
  assign n1269 = ~x96 & x125;
  assign n1270 = ~x3 & ~n1269;
  assign n1271 = ~x129 & ~n1270;
  assign n1272 = ~x126 & n713;
  assign y0 = x108;
  assign y1 = x83;
  assign y2 = x104;
  assign y3 = x103;
  assign y4 = x102;
  assign y5 = x105;
  assign y6 = x107;
  assign y7 = x101;
  assign y8 = x126;
  assign y9 = x121;
  assign y10 = x1;
  assign y11 = x0;
  assign y12 = ~1'b0;
  assign y13 = x130;
  assign y14 = x128;
  assign y15 = ~n213;
  assign y16 = n227;
  assign y17 = n259;
  assign y18 = ~n266;
  assign y19 = ~n272;
  assign y20 = ~n281;
  assign y21 = ~n285;
  assign y22 = ~n288;
  assign y23 = ~n291;
  assign y24 = ~n297;
  assign y25 = ~n300;
  assign y26 = n308;
  assign y27 = ~n312;
  assign y28 = ~n320;
  assign y29 = ~n323;
  assign y30 = n333;
  assign y31 = ~n336;
  assign y32 = ~n342;
  assign y33 = ~n347;
  assign y34 = ~n352;
  assign y35 = n372;
  assign y36 = ~n376;
  assign y37 = ~n379;
  assign y38 = n382;
  assign y39 = n398;
  assign y40 = ~n438;
  assign y41 = ~n444;
  assign y42 = n454;
  assign y43 = n466;
  assign y44 = n486;
  assign y45 = n495;
  assign y46 = n504;
  assign y47 = n513;
  assign y48 = n522;
  assign y49 = n531;
  assign y50 = n540;
  assign y51 = n549;
  assign y52 = n558;
  assign y53 = n566;
  assign y54 = n571;
  assign y55 = n579;
  assign y56 = n588;
  assign y57 = n597;
  assign y58 = n606;
  assign y59 = n612;
  assign y60 = n620;
  assign y61 = n628;
  assign y62 = n637;
  assign y63 = n646;
  assign y64 = n655;
  assign y65 = n667;
  assign y66 = n670;
  assign y67 = n673;
  assign y68 = n483;
  assign y69 = ~n674;
  assign y70 = n676;
  assign y71 = n693;
  assign y72 = n698;
  assign y73 = n701;
  assign y74 = n705;
  assign y75 = n709;
  assign y76 = n712;
  assign y77 = ~n723;
  assign y78 = ~n729;
  assign y79 = ~n735;
  assign y80 = ~n741;
  assign y81 = ~n749;
  assign y82 = ~n755;
  assign y83 = ~n761;
  assign y84 = ~n767;
  assign y85 = ~n773;
  assign y86 = ~n779;
  assign y87 = ~n785;
  assign y88 = ~n791;
  assign y89 = ~n797;
  assign y90 = ~n803;
  assign y91 = ~n809;
  assign y92 = ~n815;
  assign y93 = n823;
  assign y94 = n829;
  assign y95 = n835;
  assign y96 = n841;
  assign y97 = n847;
  assign y98 = ~n878;
  assign y99 = n884;
  assign y100 = n891;
  assign y101 = n897;
  assign y102 = n903;
  assign y103 = n911;
  assign y104 = n917;
  assign y105 = n923;
  assign y106 = n929;
  assign y107 = n935;
  assign y108 = n941;
  assign y109 = n950;
  assign y110 = n961;
  assign y111 = n970;
  assign y112 = n979;
  assign y113 = n985;
  assign y114 = n991;
  assign y115 = n1000;
  assign y116 = ~n1032;
  assign y117 = n1067;
  assign y118 = n1097;
  assign y119 = n1131;
  assign y120 = n1160;
  assign y121 = n1162;
  assign y122 = n1191;
  assign y123 = ~n1222;
  assign y124 = n1226;
  assign y125 = n1229;
  assign y126 = n1236;
  assign y127 = n1242;
  assign y128 = n1248;
  assign y129 = ~n263;
  assign y130 = n1254;
  assign y131 = n1255;
  assign y132 = ~n1256;
  assign y133 = n1259;
  assign y134 = n1260;
  assign y135 = n1263;
  assign y136 = n1265;
  assign y137 = ~n1266;
  assign y138 = ~n1267;
  assign y139 = n1268;
  assign y140 = n1271;
  assign y141 = n1272;
endmodule