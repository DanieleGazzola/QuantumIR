module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682;
  assign n129 = x0 & x64;
  assign n131 = x0 & x65;
  assign n130 = x1 & x64;
  assign n132 = n131 ^ n130;
  assign n133 = x66 ^ x2;
  assign n134 = n129 & ~n133;
  assign n135 = x2 & x64;
  assign n136 = ~x0 & ~n135;
  assign n138 = ~x64 & x66;
  assign n139 = x0 & ~n138;
  assign n137 = x1 & x65;
  assign n140 = n139 ^ n137;
  assign n141 = n140 ^ n139;
  assign n142 = ~x64 & ~x66;
  assign n143 = n142 ^ n139;
  assign n144 = ~n141 & n143;
  assign n145 = n144 ^ n139;
  assign n146 = ~n136 & ~n145;
  assign n147 = n146 ^ n137;
  assign n148 = ~n134 & n147;
  assign n165 = x64 & x65;
  assign n166 = ~x66 & ~n165;
  assign n167 = x65 & x66;
  assign n168 = ~n166 & ~n167;
  assign n169 = x2 ^ x1;
  assign n170 = ~n168 & n169;
  assign n171 = n170 ^ x1;
  assign n172 = n171 ^ x67;
  assign n158 = n133 ^ x65;
  assign n159 = n158 ^ n133;
  assign n160 = n133 ^ x66;
  assign n161 = ~n159 & n160;
  assign n162 = n161 ^ n133;
  assign n163 = ~x1 & n162;
  assign n164 = n163 ^ n133;
  assign n173 = n172 ^ n164;
  assign n174 = ~x0 & n173;
  assign n175 = n174 ^ n172;
  assign n149 = x3 & x64;
  assign n150 = n149 ^ x2;
  assign n151 = ~x0 & ~n137;
  assign n152 = ~x64 & x65;
  assign n153 = ~n138 & ~n152;
  assign n154 = ~n151 & ~n153;
  assign n155 = ~n149 & n154;
  assign n156 = n150 & n155;
  assign n157 = n156 ^ n150;
  assign n176 = n175 ^ n157;
  assign n189 = x67 & ~n166;
  assign n190 = ~x67 & ~n167;
  assign n191 = ~n189 & ~n190;
  assign n192 = n169 & ~n191;
  assign n193 = n192 ^ x1;
  assign n194 = n193 ^ x68;
  assign n187 = x67 ^ x2;
  assign n188 = x1 & n187;
  assign n195 = n194 ^ n188;
  assign n196 = n195 ^ n194;
  assign n197 = ~x1 & x2;
  assign n198 = ~x66 & n197;
  assign n199 = n198 ^ n194;
  assign n200 = n199 ^ n194;
  assign n201 = ~n196 & ~n200;
  assign n202 = n201 ^ n194;
  assign n203 = ~x0 & ~n202;
  assign n204 = n203 ^ n194;
  assign n183 = x2 & x3;
  assign n184 = n183 ^ x4;
  assign n185 = ~x64 & n184;
  assign n178 = x3 ^ x2;
  assign n179 = x65 ^ x3;
  assign n180 = n178 & ~n179;
  assign n181 = n180 ^ x2;
  assign n182 = n181 ^ x4;
  assign n186 = n185 ^ n182;
  assign n205 = n204 ^ n186;
  assign n177 = n157 & n175;
  assign n206 = n205 ^ n177;
  assign n238 = x5 ^ x4;
  assign n239 = n178 & n238;
  assign n240 = n142 & n239;
  assign n241 = x4 & ~n178;
  assign n242 = n241 ^ n183;
  assign n243 = ~n240 & ~n242;
  assign n244 = x65 & ~n243;
  assign n245 = n183 ^ x5;
  assign n246 = n245 ^ n183;
  assign n247 = ~n178 & n246;
  assign n248 = n247 ^ n183;
  assign n249 = n238 & n248;
  assign n250 = x64 & n249;
  assign n251 = n152 & n238;
  assign n252 = x66 & n178;
  assign n253 = ~n251 & n252;
  assign n254 = ~n250 & ~n253;
  assign n255 = ~n244 & n254;
  assign n233 = ~x64 & ~x65;
  assign n231 = x4 ^ x2;
  assign n232 = x64 & n231;
  assign n234 = n233 ^ n232;
  assign n235 = ~n178 & ~n234;
  assign n236 = n235 ^ n233;
  assign n237 = x5 & ~n236;
  assign n256 = n255 ^ n237;
  assign n222 = ~x68 & ~n189;
  assign n223 = x68 & ~n190;
  assign n224 = ~n222 & ~n223;
  assign n225 = n169 & ~n224;
  assign n226 = n225 ^ x1;
  assign n227 = n226 ^ x69;
  assign n210 = x68 ^ x2;
  assign n211 = n210 ^ x1;
  assign n212 = n211 ^ n210;
  assign n213 = n212 ^ x0;
  assign n214 = n210 ^ x68;
  assign n215 = n214 ^ x67;
  assign n216 = ~x67 & ~n215;
  assign n217 = n216 ^ n210;
  assign n218 = n217 ^ x67;
  assign n219 = n213 & ~n218;
  assign n220 = n219 ^ n216;
  assign n221 = n220 ^ x67;
  assign n228 = n227 ^ n221;
  assign n229 = ~x0 & ~n228;
  assign n230 = n229 ^ n227;
  assign n257 = n256 ^ n230;
  assign n207 = n186 ^ n177;
  assign n208 = n205 & ~n207;
  assign n209 = n208 ^ n204;
  assign n258 = n257 ^ n209;
  assign n279 = x66 & n242;
  assign n280 = n178 & ~n238;
  assign n281 = x67 & n280;
  assign n282 = ~n279 & ~n281;
  assign n283 = x65 & n249;
  assign n284 = n282 & ~n283;
  assign n285 = n168 ^ x67;
  assign n286 = n239 & n285;
  assign n287 = n284 & ~n286;
  assign n288 = n287 ^ x5;
  assign n289 = x6 ^ x5;
  assign n290 = n288 & n289;
  assign n291 = x5 & n236;
  assign n292 = n255 & n291;
  assign n293 = ~x6 & n292;
  assign n294 = ~n290 & ~n293;
  assign n295 = x64 & ~n294;
  assign n296 = x64 & n289;
  assign n297 = ~n292 & ~n296;
  assign n298 = n297 ^ n292;
  assign n299 = ~n288 & n298;
  assign n300 = n299 ^ n292;
  assign n301 = ~n295 & ~n300;
  assign n263 = x69 & ~n222;
  assign n264 = ~x69 & ~n223;
  assign n265 = ~n263 & ~n264;
  assign n266 = n169 & ~n265;
  assign n267 = n266 ^ x1;
  assign n268 = n267 ^ x70;
  assign n262 = ~x68 & n197;
  assign n269 = n268 ^ n262;
  assign n270 = n269 ^ n268;
  assign n271 = x69 ^ x2;
  assign n272 = x1 & n271;
  assign n273 = n272 ^ n268;
  assign n274 = n273 ^ n268;
  assign n275 = ~n270 & ~n274;
  assign n276 = n275 ^ n268;
  assign n277 = ~x0 & ~n276;
  assign n278 = n277 ^ n268;
  assign n302 = n301 ^ n278;
  assign n259 = n230 ^ n209;
  assign n260 = n257 & n259;
  assign n261 = n260 ^ n209;
  assign n303 = n302 ^ n261;
  assign n368 = ~n288 & ~n297;
  assign n321 = n191 ^ x68;
  assign n322 = n239 & n321;
  assign n323 = x67 & n242;
  assign n324 = x66 & n249;
  assign n325 = ~n323 & ~n324;
  assign n326 = x68 & n280;
  assign n327 = n325 & ~n326;
  assign n328 = ~n322 & n327;
  assign n329 = x5 & x6;
  assign n330 = n329 ^ x65;
  assign n331 = n330 ^ n329;
  assign n332 = n329 ^ x5;
  assign n333 = ~n331 & n332;
  assign n334 = n333 ^ n329;
  assign n335 = x7 & n334;
  assign n336 = n335 ^ n329;
  assign n337 = n336 ^ x5;
  assign n338 = n337 ^ n336;
  assign n340 = ~x5 & ~x6;
  assign n341 = x65 & ~n340;
  assign n339 = x7 & x64;
  assign n342 = n341 ^ n339;
  assign n343 = n342 ^ n336;
  assign n344 = n343 ^ n336;
  assign n345 = ~n338 & n344;
  assign n346 = n345 ^ n336;
  assign n347 = ~n328 & n346;
  assign n348 = n347 ^ n336;
  assign n349 = x64 & n348;
  assign n350 = n328 ^ x6;
  assign n351 = n328 ^ x5;
  assign n352 = x65 & ~n339;
  assign n353 = n352 ^ x5;
  assign n354 = x5 & n353;
  assign n355 = n354 ^ x5;
  assign n356 = ~n351 & n355;
  assign n357 = n356 ^ n354;
  assign n358 = n357 ^ x5;
  assign n359 = n358 ^ n352;
  assign n360 = n350 & n359;
  assign n361 = ~n349 & ~n360;
  assign n362 = ~x7 & x64;
  assign n363 = n362 ^ n342;
  assign n364 = n329 & n363;
  assign n365 = n364 ^ n342;
  assign n366 = n351 & ~n365;
  assign n367 = n361 & ~n366;
  assign n369 = n368 ^ n367;
  assign n312 = ~x70 & ~n263;
  assign n313 = x70 & ~n264;
  assign n314 = ~n312 & ~n313;
  assign n315 = n169 & ~n314;
  assign n316 = n315 ^ x1;
  assign n317 = n316 ^ x71;
  assign n308 = x2 & ~x69;
  assign n307 = x70 ^ x2;
  assign n309 = n308 ^ n307;
  assign n310 = x1 & n309;
  assign n311 = n310 ^ n308;
  assign n318 = n317 ^ n311;
  assign n319 = ~x0 & n318;
  assign n320 = n319 ^ n317;
  assign n370 = n369 ^ n320;
  assign n304 = n301 ^ n261;
  assign n305 = n302 & ~n304;
  assign n306 = n305 ^ n261;
  assign n371 = n370 ^ n306;
  assign n420 = n224 ^ x69;
  assign n421 = n239 & n420;
  assign n422 = x68 & n242;
  assign n423 = x67 & n249;
  assign n424 = ~n422 & ~n423;
  assign n425 = x69 & n280;
  assign n426 = n424 & ~n425;
  assign n427 = ~n421 & n426;
  assign n428 = n427 ^ x5;
  assign n398 = x8 ^ x7;
  assign n399 = n289 & n398;
  assign n400 = n142 & n399;
  assign n401 = x7 ^ x6;
  assign n402 = ~n289 & n401;
  assign n403 = ~n400 & ~n402;
  assign n404 = x65 & ~n403;
  assign n405 = n152 & n398;
  assign n406 = x66 & n289;
  assign n407 = ~n405 & n406;
  assign n408 = ~n404 & ~n407;
  assign n409 = n340 & n362;
  assign n410 = n408 & ~n409;
  assign n394 = n329 & ~n362;
  assign n395 = ~n339 & n340;
  assign n396 = ~n233 & ~n395;
  assign n397 = ~n394 & n396;
  assign n411 = n410 ^ n397;
  assign n393 = n329 & n339;
  assign n412 = n411 ^ n393;
  assign n413 = n412 ^ n411;
  assign n414 = n411 ^ n408;
  assign n415 = n414 ^ n411;
  assign n416 = ~n413 & n415;
  assign n417 = n416 ^ n411;
  assign n418 = ~x8 & n417;
  assign n419 = n418 ^ n411;
  assign n429 = n428 ^ n419;
  assign n391 = n367 & ~n368;
  assign n392 = n391 ^ n366;
  assign n430 = n429 ^ n392;
  assign n377 = x71 ^ x70;
  assign n378 = ~n314 & n377;
  assign n379 = n169 & ~n378;
  assign n380 = n379 ^ x1;
  assign n381 = n380 ^ x72;
  assign n375 = x1 & x71;
  assign n376 = n375 ^ x2;
  assign n382 = n381 ^ n376;
  assign n383 = n382 ^ n381;
  assign n384 = x70 & n197;
  assign n385 = n384 ^ n381;
  assign n386 = n385 ^ n381;
  assign n387 = n383 & ~n386;
  assign n388 = n387 ^ n381;
  assign n389 = ~x0 & n388;
  assign n390 = n389 ^ n381;
  assign n431 = n430 ^ n390;
  assign n372 = n369 ^ n306;
  assign n373 = ~n370 & n372;
  assign n374 = n373 ^ n306;
  assign n432 = n431 ^ n374;
  assign n485 = x8 & n411;
  assign n486 = n410 & n485;
  assign n469 = x66 & n402;
  assign n470 = n289 & ~n398;
  assign n471 = x67 & n470;
  assign n472 = ~n469 & ~n471;
  assign n473 = n340 ^ n329;
  assign n474 = n340 ^ x8;
  assign n475 = n474 ^ n340;
  assign n476 = n473 & ~n475;
  assign n477 = n476 ^ n340;
  assign n478 = n398 & n477;
  assign n479 = x65 & n478;
  assign n480 = n472 & ~n479;
  assign n481 = n285 & n399;
  assign n482 = n480 & ~n481;
  assign n483 = n482 ^ x8;
  assign n467 = x9 ^ x8;
  assign n468 = x64 & n467;
  assign n484 = n483 ^ n468;
  assign n487 = n486 ^ n484;
  assign n458 = n265 ^ x70;
  assign n459 = n239 & n458;
  assign n460 = x69 & n242;
  assign n461 = x70 & n280;
  assign n462 = ~n460 & ~n461;
  assign n463 = x68 & n249;
  assign n464 = n462 & ~n463;
  assign n465 = ~n459 & n464;
  assign n466 = n465 ^ x5;
  assign n488 = n487 ^ n466;
  assign n455 = n419 ^ n392;
  assign n456 = ~n429 & n455;
  assign n457 = n456 ^ n392;
  assign n489 = n488 ^ n457;
  assign n444 = x72 ^ x2;
  assign n445 = n444 ^ x71;
  assign n446 = n445 ^ n444;
  assign n447 = n444 ^ x72;
  assign n448 = ~n446 & n447;
  assign n449 = n448 ^ n444;
  assign n450 = ~x1 & n449;
  assign n451 = n450 ^ n444;
  assign n436 = x71 & ~x72;
  assign n437 = ~n312 & n436;
  assign n438 = ~x71 & x72;
  assign n439 = ~n313 & n438;
  assign n440 = ~n437 & ~n439;
  assign n441 = n169 & n440;
  assign n442 = n441 ^ x1;
  assign n443 = n442 ^ x73;
  assign n452 = n451 ^ n443;
  assign n453 = ~x0 & n452;
  assign n454 = n453 ^ n443;
  assign n490 = n489 ^ n454;
  assign n433 = n430 ^ n374;
  assign n434 = n431 & ~n433;
  assign n435 = n434 ^ n374;
  assign n491 = n490 ^ n435;
  assign n542 = ~n468 & ~n486;
  assign n543 = ~n483 & ~n542;
  assign n537 = x65 ^ x9;
  assign n538 = n467 & ~n537;
  assign n539 = n538 ^ x8;
  assign n540 = n539 ^ x10;
  assign n534 = x8 & x9;
  assign n535 = n534 ^ x10;
  assign n536 = ~x64 & n535;
  assign n541 = n540 ^ n536;
  assign n544 = n543 ^ n541;
  assign n526 = n321 & n399;
  assign n527 = x67 & n402;
  assign n528 = x66 & n478;
  assign n529 = ~n527 & ~n528;
  assign n530 = x68 & n470;
  assign n531 = n529 & ~n530;
  assign n532 = ~n526 & n531;
  assign n533 = n532 ^ x8;
  assign n545 = n544 ^ n533;
  assign n517 = n314 ^ x71;
  assign n518 = n239 & n517;
  assign n519 = x70 & n242;
  assign n520 = x69 & n249;
  assign n521 = ~n519 & ~n520;
  assign n522 = x71 & n280;
  assign n523 = n521 & ~n522;
  assign n524 = ~n518 & n523;
  assign n525 = n524 ^ x5;
  assign n546 = n545 ^ n525;
  assign n514 = n487 ^ n457;
  assign n515 = ~n488 & n514;
  assign n516 = n515 ^ n457;
  assign n547 = n546 ^ n516;
  assign n503 = ~x72 & ~n437;
  assign n504 = x73 & n503;
  assign n505 = x72 & ~x73;
  assign n506 = ~n439 & n505;
  assign n507 = ~n504 & ~n506;
  assign n508 = n169 & n507;
  assign n509 = n508 ^ x1;
  assign n510 = n509 ^ x74;
  assign n495 = x73 ^ x2;
  assign n496 = n495 ^ x72;
  assign n497 = n496 ^ n495;
  assign n498 = n495 ^ x73;
  assign n499 = ~n497 & n498;
  assign n500 = n499 ^ n495;
  assign n501 = ~x1 & n500;
  assign n502 = n501 ^ n495;
  assign n511 = n510 ^ n502;
  assign n512 = ~x0 & n511;
  assign n513 = n512 ^ n510;
  assign n548 = n547 ^ n513;
  assign n492 = n489 ^ n435;
  assign n493 = n490 & ~n492;
  assign n494 = n493 ^ n435;
  assign n549 = n548 ^ n494;
  assign n617 = x10 ^ x8;
  assign n618 = x64 & n617;
  assign n619 = n618 ^ n233;
  assign n620 = ~n467 & ~n619;
  assign n621 = n620 ^ n233;
  assign n622 = x11 & n621;
  assign n595 = x11 ^ x10;
  assign n596 = n467 & n595;
  assign n597 = n142 & n596;
  assign n598 = ~x8 & ~x9;
  assign n599 = n598 ^ n534;
  assign n600 = ~x10 & n599;
  assign n601 = n600 ^ n598;
  assign n602 = ~n597 & ~n601;
  assign n603 = x65 & ~n602;
  assign n604 = n152 & n595;
  assign n605 = x66 & n467;
  assign n606 = ~n604 & n605;
  assign n607 = ~n603 & ~n606;
  assign n611 = ~x10 & x64;
  assign n612 = n598 & n611;
  assign n613 = n607 & ~n612;
  assign n608 = x10 & x64;
  assign n609 = n534 & n608;
  assign n610 = n607 & ~n609;
  assign n614 = n613 ^ n610;
  assign n615 = ~x11 & ~n614;
  assign n616 = n615 ^ n613;
  assign n623 = n622 ^ n616;
  assign n587 = n399 & n420;
  assign n588 = x68 & n402;
  assign n589 = x67 & n478;
  assign n590 = ~n588 & ~n589;
  assign n591 = x69 & n470;
  assign n592 = n590 & ~n591;
  assign n593 = ~n587 & n592;
  assign n594 = n593 ^ x8;
  assign n624 = n623 ^ n594;
  assign n584 = n541 ^ n533;
  assign n585 = n544 & n584;
  assign n586 = n585 ^ n543;
  assign n625 = n624 ^ n586;
  assign n575 = n378 ^ x72;
  assign n576 = n239 & n575;
  assign n577 = x71 & n242;
  assign n578 = x70 & n249;
  assign n579 = ~n577 & ~n578;
  assign n580 = x72 & n280;
  assign n581 = n579 & ~n580;
  assign n582 = ~n576 & n581;
  assign n583 = n582 ^ x5;
  assign n626 = n625 ^ n583;
  assign n572 = n545 ^ n516;
  assign n573 = ~n546 & n572;
  assign n574 = n573 ^ n516;
  assign n627 = n626 ^ n574;
  assign n554 = x73 & ~n503;
  assign n555 = ~x74 & ~n554;
  assign n556 = ~x73 & ~n506;
  assign n557 = x74 & ~n556;
  assign n558 = ~n555 & ~n557;
  assign n559 = n169 & ~n558;
  assign n560 = n559 ^ x1;
  assign n561 = n560 ^ x75;
  assign n553 = ~x73 & n197;
  assign n562 = n561 ^ n553;
  assign n563 = n562 ^ n561;
  assign n564 = x74 ^ x2;
  assign n565 = x1 & n564;
  assign n566 = n565 ^ n561;
  assign n567 = n566 ^ n561;
  assign n568 = ~n563 & ~n567;
  assign n569 = n568 ^ n561;
  assign n570 = ~x0 & ~n569;
  assign n571 = n570 ^ n561;
  assign n628 = n627 ^ n571;
  assign n550 = n547 ^ n494;
  assign n551 = n548 & ~n550;
  assign n552 = n551 ^ n494;
  assign n629 = n628 ^ n552;
  assign n684 = n399 & n458;
  assign n685 = x68 & n478;
  assign n686 = x70 & n470;
  assign n687 = ~n685 & ~n686;
  assign n688 = x69 & n402;
  assign n689 = n687 & ~n688;
  assign n690 = ~n684 & n689;
  assign n691 = n690 ^ x8;
  assign n668 = x66 & n601;
  assign n669 = n534 ^ x11;
  assign n670 = n669 ^ n534;
  assign n671 = n599 & n670;
  assign n672 = n671 ^ n534;
  assign n673 = n595 & n672;
  assign n674 = x65 & n673;
  assign n675 = ~n668 & ~n674;
  assign n676 = n467 & ~n595;
  assign n677 = x67 & n676;
  assign n678 = n675 & ~n677;
  assign n679 = n285 & n596;
  assign n680 = n678 & ~n679;
  assign n681 = n680 ^ x11;
  assign n666 = x12 ^ x11;
  assign n667 = x64 & n666;
  assign n682 = n681 ^ n667;
  assign n665 = n613 & n622;
  assign n683 = n682 ^ n665;
  assign n692 = n691 ^ n683;
  assign n662 = n623 ^ n586;
  assign n663 = n624 & n662;
  assign n664 = n663 ^ n586;
  assign n693 = n692 ^ n664;
  assign n653 = n440 ^ x73;
  assign n654 = n239 & ~n653;
  assign n655 = x72 & n242;
  assign n656 = x71 & n249;
  assign n657 = ~n655 & ~n656;
  assign n658 = x73 & n280;
  assign n659 = n657 & ~n658;
  assign n660 = ~n654 & n659;
  assign n661 = n660 ^ x5;
  assign n694 = n693 ^ n661;
  assign n650 = n625 ^ n574;
  assign n651 = ~n626 & n650;
  assign n652 = n651 ^ n574;
  assign n695 = n694 ^ n652;
  assign n641 = x75 & ~n555;
  assign n642 = ~x75 & ~n557;
  assign n643 = ~n641 & ~n642;
  assign n644 = n169 & ~n643;
  assign n645 = n644 ^ x1;
  assign n646 = n645 ^ x76;
  assign n633 = x75 ^ x2;
  assign n634 = n633 ^ x74;
  assign n635 = n634 ^ n633;
  assign n636 = n633 ^ x75;
  assign n637 = ~n635 & n636;
  assign n638 = n637 ^ n633;
  assign n639 = ~x1 & n638;
  assign n640 = n639 ^ n633;
  assign n647 = n646 ^ n640;
  assign n648 = ~x0 & n647;
  assign n649 = n648 ^ n646;
  assign n696 = n695 ^ n649;
  assign n630 = n627 ^ n552;
  assign n631 = n628 & ~n630;
  assign n632 = n631 ^ n552;
  assign n697 = n696 ^ n632;
  assign n756 = ~n665 & ~n667;
  assign n757 = ~n681 & ~n756;
  assign n749 = x65 ^ x12;
  assign n750 = n666 & ~n749;
  assign n751 = n750 ^ x11;
  assign n752 = n751 ^ x13;
  assign n753 = x64 & n752;
  assign n754 = n152 & n666;
  assign n755 = ~n753 & ~n754;
  assign n758 = n757 ^ n755;
  assign n741 = n321 & n596;
  assign n742 = x66 & n673;
  assign n743 = x67 & n601;
  assign n744 = ~n742 & ~n743;
  assign n745 = x68 & n676;
  assign n746 = n744 & ~n745;
  assign n747 = ~n741 & n746;
  assign n748 = n747 ^ x11;
  assign n759 = n758 ^ n748;
  assign n733 = n399 & n517;
  assign n734 = x69 & n478;
  assign n735 = x70 & n402;
  assign n736 = ~n734 & ~n735;
  assign n737 = x71 & n470;
  assign n738 = n736 & ~n737;
  assign n739 = ~n733 & n738;
  assign n740 = n739 ^ x8;
  assign n760 = n759 ^ n740;
  assign n730 = n691 ^ n664;
  assign n731 = ~n692 & ~n730;
  assign n732 = n731 ^ n664;
  assign n761 = n760 ^ n732;
  assign n721 = n507 ^ x74;
  assign n722 = n239 & ~n721;
  assign n723 = x73 & n242;
  assign n724 = x74 & n280;
  assign n725 = ~n723 & ~n724;
  assign n726 = x72 & n249;
  assign n727 = n725 & ~n726;
  assign n728 = ~n722 & n727;
  assign n729 = n728 ^ x5;
  assign n762 = n761 ^ n729;
  assign n718 = n693 ^ n652;
  assign n719 = n694 & ~n718;
  assign n720 = n719 ^ n652;
  assign n763 = n762 ^ n720;
  assign n703 = ~x76 & ~n641;
  assign n704 = x76 & ~n642;
  assign n705 = ~n703 & ~n704;
  assign n706 = n169 & ~n705;
  assign n707 = n706 ^ x1;
  assign n708 = n707 ^ x77;
  assign n701 = x76 ^ x2;
  assign n702 = x1 & n701;
  assign n709 = n708 ^ n702;
  assign n710 = n709 ^ n708;
  assign n711 = ~x75 & n197;
  assign n712 = n711 ^ n708;
  assign n713 = n712 ^ n708;
  assign n714 = ~n710 & ~n713;
  assign n715 = n714 ^ n708;
  assign n716 = ~x0 & ~n715;
  assign n717 = n716 ^ n708;
  assign n764 = n763 ^ n717;
  assign n698 = n695 ^ n632;
  assign n699 = ~n696 & n698;
  assign n700 = n699 ^ n632;
  assign n765 = n764 ^ n700;
  assign n832 = n420 & n596;
  assign n833 = x67 & n673;
  assign n834 = x68 & n601;
  assign n835 = ~n833 & ~n834;
  assign n836 = x69 & n676;
  assign n837 = n835 & ~n836;
  assign n838 = ~n832 & n837;
  assign n839 = n838 ^ x11;
  assign n820 = x14 ^ x13;
  assign n821 = n666 & n820;
  assign n822 = n142 & n821;
  assign n823 = x13 & ~n666;
  assign n813 = x11 & x12;
  assign n824 = n823 ^ n813;
  assign n825 = ~n822 & ~n824;
  assign n826 = x65 & ~n825;
  assign n827 = n152 & n820;
  assign n828 = x66 & n666;
  assign n829 = ~n827 & n828;
  assign n830 = ~n826 & ~n829;
  assign n812 = ~x64 & ~n754;
  assign n814 = x13 & x64;
  assign n815 = n813 & n814;
  assign n816 = ~n812 & ~n815;
  assign n817 = n816 ^ n815;
  assign n818 = x14 & n817;
  assign n819 = n818 ^ n815;
  assign n831 = n830 ^ n819;
  assign n840 = n839 ^ n831;
  assign n809 = n755 ^ n748;
  assign n810 = ~n758 & ~n809;
  assign n811 = n810 ^ n757;
  assign n841 = n840 ^ n811;
  assign n801 = n399 & n575;
  assign n802 = x71 & n402;
  assign n803 = x70 & n478;
  assign n804 = ~n802 & ~n803;
  assign n805 = x72 & n470;
  assign n806 = n804 & ~n805;
  assign n807 = ~n801 & n806;
  assign n808 = n807 ^ x8;
  assign n842 = n841 ^ n808;
  assign n798 = n759 ^ n732;
  assign n799 = n760 & n798;
  assign n800 = n799 ^ n732;
  assign n843 = n842 ^ n800;
  assign n789 = n558 ^ x75;
  assign n790 = n239 & n789;
  assign n791 = x73 & n249;
  assign n792 = x74 & n242;
  assign n793 = ~n791 & ~n792;
  assign n794 = x75 & n280;
  assign n795 = n793 & ~n794;
  assign n796 = ~n790 & n795;
  assign n797 = n796 ^ x5;
  assign n844 = n843 ^ n797;
  assign n786 = n761 ^ n720;
  assign n787 = ~n762 & n786;
  assign n788 = n787 ^ n720;
  assign n845 = n844 ^ n788;
  assign n770 = x77 & ~n703;
  assign n771 = ~x77 & ~n704;
  assign n772 = ~n770 & ~n771;
  assign n773 = n169 & ~n772;
  assign n774 = n773 ^ x1;
  assign n775 = n774 ^ x78;
  assign n769 = ~x76 & n197;
  assign n776 = n775 ^ n769;
  assign n777 = n776 ^ n775;
  assign n778 = x77 ^ x2;
  assign n779 = x1 & n778;
  assign n780 = n779 ^ n775;
  assign n781 = n780 ^ n775;
  assign n782 = ~n777 & ~n781;
  assign n783 = n782 ^ n775;
  assign n784 = ~x0 & ~n783;
  assign n785 = n784 ^ n775;
  assign n846 = n845 ^ n785;
  assign n766 = n763 ^ n700;
  assign n767 = n764 & ~n766;
  assign n768 = n767 ^ n700;
  assign n847 = n846 ^ n768;
  assign n913 = n458 & n596;
  assign n914 = x69 & n601;
  assign n915 = x68 & n673;
  assign n916 = ~n914 & ~n915;
  assign n917 = x70 & n676;
  assign n918 = n916 & ~n917;
  assign n919 = ~n913 & n918;
  assign n920 = n919 ^ x11;
  assign n909 = x14 & ~n816;
  assign n910 = n830 & n909;
  assign n907 = x15 ^ x14;
  assign n908 = x64 & n907;
  assign n911 = n910 ^ n908;
  assign n893 = x66 & n824;
  assign n894 = n813 ^ x14;
  assign n895 = n894 ^ n813;
  assign n896 = ~n666 & n895;
  assign n897 = n896 ^ n813;
  assign n898 = n820 & n897;
  assign n899 = x65 & n898;
  assign n900 = ~n893 & ~n899;
  assign n901 = n666 & ~n820;
  assign n902 = x67 & n901;
  assign n903 = n900 & ~n902;
  assign n904 = n285 & n821;
  assign n905 = n903 & ~n904;
  assign n906 = n905 ^ x14;
  assign n912 = n911 ^ n906;
  assign n921 = n920 ^ n912;
  assign n890 = n839 ^ n811;
  assign n891 = ~n840 & ~n890;
  assign n892 = n891 ^ n811;
  assign n922 = n921 ^ n892;
  assign n882 = n399 & ~n653;
  assign n883 = x72 & n402;
  assign n884 = x71 & n478;
  assign n885 = ~n883 & ~n884;
  assign n886 = x73 & n470;
  assign n887 = n885 & ~n886;
  assign n888 = ~n882 & n887;
  assign n889 = n888 ^ x8;
  assign n923 = n922 ^ n889;
  assign n879 = n841 ^ n800;
  assign n880 = n842 & n879;
  assign n881 = n880 ^ n800;
  assign n924 = n923 ^ n881;
  assign n870 = n643 ^ x76;
  assign n871 = n239 & n870;
  assign n872 = x74 & n249;
  assign n873 = x75 & n242;
  assign n874 = ~n872 & ~n873;
  assign n875 = x76 & n280;
  assign n876 = n874 & ~n875;
  assign n877 = ~n871 & n876;
  assign n878 = n877 ^ x5;
  assign n925 = n924 ^ n878;
  assign n867 = n843 ^ n788;
  assign n868 = ~n844 & n867;
  assign n869 = n868 ^ n788;
  assign n926 = n925 ^ n869;
  assign n859 = x78 ^ x77;
  assign n860 = ~n772 & n859;
  assign n861 = n169 & ~n860;
  assign n862 = n861 ^ x1;
  assign n863 = n862 ^ x79;
  assign n851 = x78 ^ x2;
  assign n852 = n851 ^ x77;
  assign n853 = n852 ^ n851;
  assign n854 = n851 ^ x78;
  assign n855 = ~n853 & n854;
  assign n856 = n855 ^ n851;
  assign n857 = ~x1 & n856;
  assign n858 = n857 ^ n851;
  assign n864 = n863 ^ n858;
  assign n865 = ~x0 & n864;
  assign n866 = n865 ^ n863;
  assign n927 = n926 ^ n866;
  assign n848 = n845 ^ n768;
  assign n849 = n846 & ~n848;
  assign n850 = n849 ^ n768;
  assign n928 = n927 ^ n850;
  assign n1001 = x14 & x15;
  assign n1002 = n1001 ^ x16;
  assign n1003 = ~x64 & n1002;
  assign n997 = x65 ^ x15;
  assign n998 = n907 & ~n997;
  assign n999 = n998 ^ x14;
  assign n1000 = n999 ^ x16;
  assign n1004 = n1003 ^ n1000;
  assign n995 = ~n908 & ~n910;
  assign n996 = ~n906 & ~n995;
  assign n1005 = n1004 ^ n996;
  assign n987 = n321 & n821;
  assign n988 = x67 & n824;
  assign n989 = x66 & n898;
  assign n990 = ~n988 & ~n989;
  assign n991 = x68 & n901;
  assign n992 = n990 & ~n991;
  assign n993 = ~n987 & n992;
  assign n994 = n993 ^ x14;
  assign n1006 = n1005 ^ n994;
  assign n979 = n517 & n596;
  assign n980 = x69 & n673;
  assign n981 = x70 & n601;
  assign n982 = ~n980 & ~n981;
  assign n983 = x71 & n676;
  assign n984 = n982 & ~n983;
  assign n985 = ~n979 & n984;
  assign n986 = n985 ^ x11;
  assign n1007 = n1006 ^ n986;
  assign n976 = n920 ^ n892;
  assign n977 = ~n921 & ~n976;
  assign n978 = n977 ^ n892;
  assign n1008 = n1007 ^ n978;
  assign n968 = n399 & ~n721;
  assign n969 = x73 & n402;
  assign n970 = x72 & n478;
  assign n971 = ~n969 & ~n970;
  assign n972 = x74 & n470;
  assign n973 = n971 & ~n972;
  assign n974 = ~n968 & n973;
  assign n975 = n974 ^ x8;
  assign n1009 = n1008 ^ n975;
  assign n965 = n922 ^ n881;
  assign n966 = n923 & n965;
  assign n967 = n966 ^ n881;
  assign n1010 = n1009 ^ n967;
  assign n956 = n705 ^ x77;
  assign n957 = n239 & n956;
  assign n958 = x75 & n249;
  assign n959 = x76 & n242;
  assign n960 = ~n958 & ~n959;
  assign n961 = x77 & n280;
  assign n962 = n960 & ~n961;
  assign n963 = ~n957 & n962;
  assign n964 = n963 ^ x5;
  assign n1011 = n1010 ^ n964;
  assign n953 = n924 ^ n869;
  assign n954 = ~n925 & n953;
  assign n955 = n954 ^ n869;
  assign n1012 = n1011 ^ n955;
  assign n934 = x79 ^ x78;
  assign n935 = n771 ^ n770;
  assign n936 = n770 ^ x79;
  assign n937 = n936 ^ n770;
  assign n938 = n935 & ~n937;
  assign n939 = n938 ^ n770;
  assign n940 = n934 & ~n939;
  assign n941 = n169 & ~n940;
  assign n942 = n941 ^ x1;
  assign n943 = n942 ^ x80;
  assign n932 = x79 ^ x2;
  assign n933 = x1 & n932;
  assign n944 = n943 ^ n933;
  assign n945 = n944 ^ n943;
  assign n946 = ~x78 & n197;
  assign n947 = n946 ^ n943;
  assign n948 = n947 ^ n943;
  assign n949 = ~n945 & ~n948;
  assign n950 = n949 ^ n943;
  assign n951 = ~x0 & ~n950;
  assign n952 = n951 ^ n943;
  assign n1013 = n1012 ^ n952;
  assign n929 = n926 ^ n850;
  assign n930 = n927 & ~n929;
  assign n931 = n930 ^ n850;
  assign n1014 = n1013 ^ n931;
  assign n1083 = ~x14 & ~x15;
  assign n1094 = ~x16 & x17;
  assign n1095 = n1083 & n1094;
  assign n1096 = x64 & n1095;
  assign n1097 = x17 ^ x16;
  assign n1098 = n907 & n1097;
  assign n1099 = n142 & n1098;
  assign n1100 = n1083 ^ n1001;
  assign n1101 = x16 & n1100;
  assign n1102 = n1101 ^ n1001;
  assign n1103 = ~n1099 & ~n1102;
  assign n1104 = x65 & ~n1103;
  assign n1105 = n152 & n1097;
  assign n1106 = x66 & n907;
  assign n1107 = ~n1105 & n1106;
  assign n1108 = ~n1104 & ~n1107;
  assign n1109 = n1108 ^ x17;
  assign n1110 = x16 & x64;
  assign n1111 = n1001 & n1110;
  assign n1112 = n1108 & n1111;
  assign n1113 = n1109 & n1112;
  assign n1114 = n1113 ^ n1109;
  assign n1115 = ~n1096 & ~n1114;
  assign n1084 = ~n233 & ~n1083;
  assign n1085 = n1084 ^ n1001;
  assign n1086 = x64 ^ x16;
  assign n1087 = n1086 ^ x16;
  assign n1088 = n1084 ^ x16;
  assign n1089 = ~n1087 & n1088;
  assign n1090 = n1089 ^ x16;
  assign n1091 = ~n1085 & ~n1090;
  assign n1092 = n1091 ^ n1001;
  assign n1093 = x17 & n1092;
  assign n1116 = n1115 ^ n1093;
  assign n1075 = n420 & n821;
  assign n1076 = x68 & n824;
  assign n1077 = x67 & n898;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = x69 & n901;
  assign n1080 = n1078 & ~n1079;
  assign n1081 = ~n1075 & n1080;
  assign n1082 = n1081 ^ x14;
  assign n1117 = n1116 ^ n1082;
  assign n1072 = n1004 ^ n994;
  assign n1073 = n1005 & n1072;
  assign n1074 = n1073 ^ n996;
  assign n1118 = n1117 ^ n1074;
  assign n1064 = n575 & n596;
  assign n1065 = x71 & n601;
  assign n1066 = x70 & n673;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = x72 & n676;
  assign n1069 = n1067 & ~n1068;
  assign n1070 = ~n1064 & n1069;
  assign n1071 = n1070 ^ x11;
  assign n1119 = n1118 ^ n1071;
  assign n1061 = n1006 ^ n978;
  assign n1062 = ~n1007 & ~n1061;
  assign n1063 = n1062 ^ n978;
  assign n1120 = n1119 ^ n1063;
  assign n1053 = n399 & n789;
  assign n1054 = x74 & n402;
  assign n1055 = x73 & n478;
  assign n1056 = ~n1054 & ~n1055;
  assign n1057 = x75 & n470;
  assign n1058 = n1056 & ~n1057;
  assign n1059 = ~n1053 & n1058;
  assign n1060 = n1059 ^ x8;
  assign n1121 = n1120 ^ n1060;
  assign n1050 = n1008 ^ n967;
  assign n1051 = n1009 & n1050;
  assign n1052 = n1051 ^ n967;
  assign n1122 = n1121 ^ n1052;
  assign n1041 = n772 ^ x78;
  assign n1042 = n239 & n1041;
  assign n1043 = x76 & n249;
  assign n1044 = x78 & n280;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = x77 & n242;
  assign n1047 = n1045 & ~n1046;
  assign n1048 = ~n1042 & n1047;
  assign n1049 = n1048 ^ x5;
  assign n1123 = n1122 ^ n1049;
  assign n1038 = n1010 ^ n955;
  assign n1039 = ~n1011 & n1038;
  assign n1040 = n1039 ^ n955;
  assign n1124 = n1123 ^ n1040;
  assign n1030 = x80 ^ x79;
  assign n1031 = ~n940 & n1030;
  assign n1032 = n169 & ~n1031;
  assign n1033 = n1032 ^ x1;
  assign n1034 = n1033 ^ x81;
  assign n1018 = x80 ^ x2;
  assign n1019 = n1018 ^ x1;
  assign n1020 = n1019 ^ n1018;
  assign n1021 = n1020 ^ x0;
  assign n1022 = n1018 ^ x80;
  assign n1023 = n1022 ^ x79;
  assign n1024 = ~x79 & ~n1023;
  assign n1025 = n1024 ^ n1018;
  assign n1026 = n1025 ^ x79;
  assign n1027 = n1021 & ~n1026;
  assign n1028 = n1027 ^ n1024;
  assign n1029 = n1028 ^ x79;
  assign n1035 = n1034 ^ n1029;
  assign n1036 = ~x0 & ~n1035;
  assign n1037 = n1036 ^ n1034;
  assign n1125 = n1124 ^ n1037;
  assign n1015 = n1012 ^ n931;
  assign n1016 = n1013 & ~n1015;
  assign n1017 = n1016 ^ n931;
  assign n1126 = n1125 ^ n1017;
  assign n1208 = n1093 & n1115;
  assign n1193 = x66 & n1102;
  assign n1194 = n1001 ^ x17;
  assign n1195 = n1194 ^ n1001;
  assign n1196 = n1100 & n1195;
  assign n1197 = n1196 ^ n1001;
  assign n1198 = n1097 & n1197;
  assign n1199 = x65 & n1198;
  assign n1200 = ~n1193 & ~n1199;
  assign n1201 = n907 & ~n1097;
  assign n1202 = x67 & n1201;
  assign n1203 = n1200 & ~n1202;
  assign n1204 = n285 & n1098;
  assign n1205 = n1203 & ~n1204;
  assign n1206 = n1205 ^ x17;
  assign n1191 = x18 ^ x17;
  assign n1192 = x64 & n1191;
  assign n1207 = n1206 ^ n1192;
  assign n1209 = n1208 ^ n1207;
  assign n1183 = n458 & n821;
  assign n1184 = x69 & n824;
  assign n1185 = x68 & n898;
  assign n1186 = ~n1184 & ~n1185;
  assign n1187 = x70 & n901;
  assign n1188 = n1186 & ~n1187;
  assign n1189 = ~n1183 & n1188;
  assign n1190 = n1189 ^ x14;
  assign n1210 = n1209 ^ n1190;
  assign n1180 = n1116 ^ n1074;
  assign n1181 = n1117 & n1180;
  assign n1182 = n1181 ^ n1074;
  assign n1211 = n1210 ^ n1182;
  assign n1172 = n596 & ~n653;
  assign n1173 = x71 & n673;
  assign n1174 = x73 & n676;
  assign n1175 = ~n1173 & ~n1174;
  assign n1176 = x72 & n601;
  assign n1177 = n1175 & ~n1176;
  assign n1178 = ~n1172 & n1177;
  assign n1179 = n1178 ^ x11;
  assign n1212 = n1211 ^ n1179;
  assign n1169 = n1118 ^ n1063;
  assign n1170 = ~n1119 & ~n1169;
  assign n1171 = n1170 ^ n1063;
  assign n1213 = n1212 ^ n1171;
  assign n1161 = n399 & n870;
  assign n1162 = x74 & n478;
  assign n1163 = x75 & n402;
  assign n1164 = ~n1162 & ~n1163;
  assign n1165 = x76 & n470;
  assign n1166 = n1164 & ~n1165;
  assign n1167 = ~n1161 & n1166;
  assign n1168 = n1167 ^ x8;
  assign n1214 = n1213 ^ n1168;
  assign n1158 = n1120 ^ n1052;
  assign n1159 = n1121 & n1158;
  assign n1160 = n1159 ^ n1052;
  assign n1215 = n1214 ^ n1160;
  assign n1149 = n860 ^ x79;
  assign n1150 = n239 & n1149;
  assign n1151 = x77 & n249;
  assign n1152 = x79 & n280;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = x78 & n242;
  assign n1155 = n1153 & ~n1154;
  assign n1156 = ~n1150 & n1155;
  assign n1157 = n1156 ^ x5;
  assign n1216 = n1215 ^ n1157;
  assign n1146 = n1122 ^ n1040;
  assign n1147 = ~n1123 & n1146;
  assign n1148 = n1147 ^ n1040;
  assign n1217 = n1216 ^ n1148;
  assign n1135 = x81 ^ x2;
  assign n1136 = n1135 ^ x81;
  assign n1137 = n1135 ^ x80;
  assign n1138 = n1137 ^ n1135;
  assign n1139 = n1136 & ~n1138;
  assign n1140 = n1139 ^ n1135;
  assign n1141 = ~x1 & n1140;
  assign n1142 = n1141 ^ n1135;
  assign n1130 = x81 ^ x80;
  assign n1131 = ~n1031 & n1130;
  assign n1132 = n169 & ~n1131;
  assign n1133 = n1132 ^ x1;
  assign n1134 = n1133 ^ x82;
  assign n1143 = n1142 ^ n1134;
  assign n1144 = ~x0 & n1143;
  assign n1145 = n1144 ^ n1134;
  assign n1218 = n1217 ^ n1145;
  assign n1127 = n1124 ^ n1017;
  assign n1128 = n1125 & ~n1127;
  assign n1129 = n1128 ^ n1017;
  assign n1219 = n1218 ^ n1129;
  assign n1301 = ~n1192 & ~n1208;
  assign n1302 = ~n1206 & ~n1301;
  assign n1292 = n321 & n1098;
  assign n1293 = x67 & n1102;
  assign n1294 = x66 & n1198;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = x68 & n1201;
  assign n1297 = n1295 & ~n1296;
  assign n1298 = ~n1292 & n1297;
  assign n1299 = n1298 ^ x17;
  assign n1287 = x65 ^ x18;
  assign n1288 = n1191 & ~n1287;
  assign n1289 = n1288 ^ x17;
  assign n1290 = n1289 ^ x19;
  assign n1284 = x17 & x18;
  assign n1285 = n1284 ^ x19;
  assign n1286 = ~x64 & n1285;
  assign n1291 = n1290 ^ n1286;
  assign n1300 = n1299 ^ n1291;
  assign n1303 = n1302 ^ n1300;
  assign n1276 = n517 & n821;
  assign n1277 = x70 & n824;
  assign n1278 = x69 & n898;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = x71 & n901;
  assign n1281 = n1279 & ~n1280;
  assign n1282 = ~n1276 & n1281;
  assign n1283 = n1282 ^ x14;
  assign n1304 = n1303 ^ n1283;
  assign n1273 = n1209 ^ n1182;
  assign n1274 = ~n1210 & ~n1273;
  assign n1275 = n1274 ^ n1182;
  assign n1305 = n1304 ^ n1275;
  assign n1265 = n596 & ~n721;
  assign n1266 = x73 & n601;
  assign n1267 = x72 & n673;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = x74 & n676;
  assign n1270 = n1268 & ~n1269;
  assign n1271 = ~n1265 & n1270;
  assign n1272 = n1271 ^ x11;
  assign n1306 = n1305 ^ n1272;
  assign n1262 = n1211 ^ n1171;
  assign n1263 = n1212 & n1262;
  assign n1264 = n1263 ^ n1171;
  assign n1307 = n1306 ^ n1264;
  assign n1254 = n399 & n956;
  assign n1255 = x75 & n478;
  assign n1256 = x76 & n402;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = x77 & n470;
  assign n1259 = n1257 & ~n1258;
  assign n1260 = ~n1254 & n1259;
  assign n1261 = n1260 ^ x8;
  assign n1308 = n1307 ^ n1261;
  assign n1251 = n1213 ^ n1160;
  assign n1252 = ~n1214 & ~n1251;
  assign n1253 = n1252 ^ n1160;
  assign n1309 = n1308 ^ n1253;
  assign n1242 = n940 ^ x80;
  assign n1243 = n239 & n1242;
  assign n1244 = x79 & n242;
  assign n1245 = x80 & n280;
  assign n1246 = ~n1244 & ~n1245;
  assign n1247 = x78 & n249;
  assign n1248 = n1246 & ~n1247;
  assign n1249 = ~n1243 & n1248;
  assign n1250 = n1249 ^ x5;
  assign n1310 = n1309 ^ n1250;
  assign n1239 = n1215 ^ n1148;
  assign n1240 = n1216 & ~n1239;
  assign n1241 = n1240 ^ n1148;
  assign n1311 = n1310 ^ n1241;
  assign n1225 = x82 ^ x81;
  assign n1226 = ~n1131 & n1225;
  assign n1227 = n169 & ~n1226;
  assign n1228 = n1227 ^ x1;
  assign n1229 = n1228 ^ x83;
  assign n1223 = x82 ^ x2;
  assign n1224 = x1 & n1223;
  assign n1230 = n1229 ^ n1224;
  assign n1231 = n1230 ^ n1229;
  assign n1232 = ~x81 & n197;
  assign n1233 = n1232 ^ n1229;
  assign n1234 = n1233 ^ n1229;
  assign n1235 = ~n1231 & ~n1234;
  assign n1236 = n1235 ^ n1229;
  assign n1237 = ~x0 & ~n1236;
  assign n1238 = n1237 ^ n1229;
  assign n1312 = n1311 ^ n1238;
  assign n1220 = n1217 ^ n1129;
  assign n1221 = ~n1218 & n1220;
  assign n1222 = n1221 ^ n1129;
  assign n1313 = n1312 ^ n1222;
  assign n1399 = ~x17 & ~x18;
  assign n1400 = ~x19 & x20;
  assign n1401 = n1399 & n1400;
  assign n1402 = x64 & n1401;
  assign n1403 = x20 ^ x19;
  assign n1404 = n1191 & n1403;
  assign n1405 = n142 & n1404;
  assign n1406 = n1399 ^ n1284;
  assign n1407 = x19 & n1406;
  assign n1408 = n1407 ^ n1284;
  assign n1409 = ~n1405 & ~n1408;
  assign n1410 = x65 & ~n1409;
  assign n1411 = n152 & n1403;
  assign n1412 = x66 & n1191;
  assign n1413 = ~n1411 & n1412;
  assign n1414 = ~n1410 & ~n1413;
  assign n1415 = n1414 ^ x20;
  assign n1416 = x19 & x64;
  assign n1417 = n1284 & n1416;
  assign n1418 = n1414 & n1417;
  assign n1419 = n1415 & n1418;
  assign n1420 = n1419 ^ n1415;
  assign n1421 = ~n1402 & ~n1420;
  assign n1393 = x19 ^ x17;
  assign n1394 = x64 & n1393;
  assign n1395 = n1394 ^ n233;
  assign n1396 = ~n1191 & ~n1395;
  assign n1397 = n1396 ^ n233;
  assign n1398 = x20 & n1397;
  assign n1422 = n1421 ^ n1398;
  assign n1385 = n420 & n1098;
  assign n1386 = x67 & n1198;
  assign n1387 = x69 & n1201;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = x68 & n1102;
  assign n1390 = n1388 & ~n1389;
  assign n1391 = ~n1385 & n1390;
  assign n1392 = n1391 ^ x17;
  assign n1423 = n1422 ^ n1392;
  assign n1382 = n1302 ^ n1299;
  assign n1383 = n1300 & ~n1382;
  assign n1384 = n1383 ^ n1302;
  assign n1424 = n1423 ^ n1384;
  assign n1374 = n575 & n821;
  assign n1375 = x71 & n824;
  assign n1376 = x70 & n898;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = x72 & n901;
  assign n1379 = n1377 & ~n1378;
  assign n1380 = ~n1374 & n1379;
  assign n1381 = n1380 ^ x14;
  assign n1425 = n1424 ^ n1381;
  assign n1371 = n1303 ^ n1275;
  assign n1372 = ~n1304 & ~n1371;
  assign n1373 = n1372 ^ n1275;
  assign n1426 = n1425 ^ n1373;
  assign n1363 = n596 & n789;
  assign n1364 = x73 & n673;
  assign n1365 = x75 & n676;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = x74 & n601;
  assign n1368 = n1366 & ~n1367;
  assign n1369 = ~n1363 & n1368;
  assign n1370 = n1369 ^ x11;
  assign n1427 = n1426 ^ n1370;
  assign n1360 = n1305 ^ n1264;
  assign n1361 = n1306 & n1360;
  assign n1362 = n1361 ^ n1264;
  assign n1428 = n1427 ^ n1362;
  assign n1352 = n399 & n1041;
  assign n1353 = x76 & n478;
  assign n1354 = x78 & n470;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = x77 & n402;
  assign n1357 = n1355 & ~n1356;
  assign n1358 = ~n1352 & n1357;
  assign n1359 = n1358 ^ x8;
  assign n1429 = n1428 ^ n1359;
  assign n1349 = n1307 ^ n1253;
  assign n1350 = ~n1308 & ~n1349;
  assign n1351 = n1350 ^ n1253;
  assign n1430 = n1429 ^ n1351;
  assign n1340 = n1031 ^ x81;
  assign n1341 = n239 & n1340;
  assign n1342 = x79 & n249;
  assign n1343 = x80 & n242;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = x81 & n280;
  assign n1346 = n1344 & ~n1345;
  assign n1347 = ~n1341 & n1346;
  assign n1348 = n1347 ^ x5;
  assign n1431 = n1430 ^ n1348;
  assign n1337 = n1309 ^ n1241;
  assign n1338 = n1310 & ~n1337;
  assign n1339 = n1338 ^ n1241;
  assign n1432 = n1431 ^ n1339;
  assign n1329 = x83 ^ x82;
  assign n1330 = ~n1226 & n1329;
  assign n1331 = n169 & ~n1330;
  assign n1332 = n1331 ^ x1;
  assign n1333 = n1332 ^ x84;
  assign n1317 = x83 ^ x2;
  assign n1318 = n1317 ^ x1;
  assign n1319 = n1318 ^ n1317;
  assign n1320 = n1319 ^ x0;
  assign n1321 = n1317 ^ x83;
  assign n1322 = n1321 ^ x82;
  assign n1323 = ~x82 & ~n1322;
  assign n1324 = n1323 ^ n1317;
  assign n1325 = n1324 ^ x82;
  assign n1326 = n1320 & ~n1325;
  assign n1327 = n1326 ^ n1323;
  assign n1328 = n1327 ^ x82;
  assign n1334 = n1333 ^ n1328;
  assign n1335 = ~x0 & ~n1334;
  assign n1336 = n1335 ^ n1333;
  assign n1433 = n1432 ^ n1336;
  assign n1314 = n1311 ^ n1222;
  assign n1315 = ~n1312 & n1314;
  assign n1316 = n1315 ^ n1222;
  assign n1434 = n1433 ^ n1316;
  assign n1524 = n1398 & n1421;
  assign n1509 = x66 & n1408;
  assign n1510 = n1284 ^ x20;
  assign n1511 = n1510 ^ n1284;
  assign n1512 = n1406 & n1511;
  assign n1513 = n1512 ^ n1284;
  assign n1514 = n1403 & n1513;
  assign n1515 = x65 & n1514;
  assign n1516 = ~n1509 & ~n1515;
  assign n1517 = n1191 & ~n1403;
  assign n1518 = x67 & n1517;
  assign n1519 = n1516 & ~n1518;
  assign n1520 = n285 & n1404;
  assign n1521 = n1519 & ~n1520;
  assign n1522 = n1521 ^ x20;
  assign n1507 = x21 ^ x20;
  assign n1508 = x64 & n1507;
  assign n1523 = n1522 ^ n1508;
  assign n1525 = n1524 ^ n1523;
  assign n1499 = n458 & n1098;
  assign n1500 = x68 & n1198;
  assign n1501 = x70 & n1201;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = x69 & n1102;
  assign n1504 = n1502 & ~n1503;
  assign n1505 = ~n1499 & n1504;
  assign n1506 = n1505 ^ x17;
  assign n1526 = n1525 ^ n1506;
  assign n1496 = n1422 ^ n1384;
  assign n1497 = n1423 & n1496;
  assign n1498 = n1497 ^ n1384;
  assign n1527 = n1526 ^ n1498;
  assign n1488 = ~n653 & n821;
  assign n1489 = x71 & n898;
  assign n1490 = x73 & n901;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = x72 & n824;
  assign n1493 = n1491 & ~n1492;
  assign n1494 = ~n1488 & n1493;
  assign n1495 = n1494 ^ x14;
  assign n1528 = n1527 ^ n1495;
  assign n1485 = n1424 ^ n1373;
  assign n1486 = ~n1425 & ~n1485;
  assign n1487 = n1486 ^ n1373;
  assign n1529 = n1528 ^ n1487;
  assign n1477 = n596 & n870;
  assign n1478 = x75 & n601;
  assign n1479 = x76 & n676;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = x74 & n673;
  assign n1482 = n1480 & ~n1481;
  assign n1483 = ~n1477 & n1482;
  assign n1484 = n1483 ^ x11;
  assign n1530 = n1529 ^ n1484;
  assign n1474 = n1426 ^ n1362;
  assign n1475 = n1427 & n1474;
  assign n1476 = n1475 ^ n1362;
  assign n1531 = n1530 ^ n1476;
  assign n1466 = n399 & n1149;
  assign n1467 = x77 & n478;
  assign n1468 = x78 & n402;
  assign n1469 = ~n1467 & ~n1468;
  assign n1470 = x79 & n470;
  assign n1471 = n1469 & ~n1470;
  assign n1472 = ~n1466 & n1471;
  assign n1473 = n1472 ^ x8;
  assign n1532 = n1531 ^ n1473;
  assign n1463 = n1428 ^ n1351;
  assign n1464 = ~n1429 & ~n1463;
  assign n1465 = n1464 ^ n1351;
  assign n1533 = n1532 ^ n1465;
  assign n1454 = n1131 ^ x82;
  assign n1455 = n239 & n1454;
  assign n1456 = x80 & n249;
  assign n1457 = x81 & n242;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = x82 & n280;
  assign n1460 = n1458 & ~n1459;
  assign n1461 = ~n1455 & n1460;
  assign n1462 = n1461 ^ x5;
  assign n1534 = n1533 ^ n1462;
  assign n1451 = n1430 ^ n1339;
  assign n1452 = n1431 & ~n1451;
  assign n1453 = n1452 ^ n1339;
  assign n1535 = n1534 ^ n1453;
  assign n1443 = x84 ^ x83;
  assign n1444 = ~n1330 & n1443;
  assign n1445 = n169 & ~n1444;
  assign n1446 = n1445 ^ x1;
  assign n1447 = n1446 ^ x85;
  assign n1439 = x2 & ~x83;
  assign n1438 = x84 ^ x2;
  assign n1440 = n1439 ^ n1438;
  assign n1441 = x1 & n1440;
  assign n1442 = n1441 ^ n1439;
  assign n1448 = n1447 ^ n1442;
  assign n1449 = ~x0 & n1448;
  assign n1450 = n1449 ^ n1447;
  assign n1536 = n1535 ^ n1450;
  assign n1435 = n1432 ^ n1316;
  assign n1436 = ~n1433 & n1435;
  assign n1437 = n1436 ^ n1316;
  assign n1537 = n1536 ^ n1437;
  assign n1630 = ~n1508 & ~n1524;
  assign n1631 = ~n1522 & ~n1630;
  assign n1625 = x20 & x21;
  assign n1626 = n1625 ^ x22;
  assign n1627 = ~x64 & n1626;
  assign n1621 = x65 ^ x21;
  assign n1622 = n1507 & ~n1621;
  assign n1623 = n1622 ^ x20;
  assign n1624 = n1623 ^ x22;
  assign n1628 = n1627 ^ n1624;
  assign n1613 = n321 & n1404;
  assign n1614 = x66 & n1514;
  assign n1615 = x68 & n1517;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = x67 & n1408;
  assign n1618 = n1616 & ~n1617;
  assign n1619 = ~n1613 & n1618;
  assign n1620 = n1619 ^ x20;
  assign n1629 = n1628 ^ n1620;
  assign n1632 = n1631 ^ n1629;
  assign n1605 = n517 & n1098;
  assign n1606 = x69 & n1198;
  assign n1607 = x71 & n1201;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = x70 & n1102;
  assign n1610 = n1608 & ~n1609;
  assign n1611 = ~n1605 & n1610;
  assign n1612 = n1611 ^ x17;
  assign n1633 = n1632 ^ n1612;
  assign n1602 = n1525 ^ n1498;
  assign n1603 = ~n1526 & ~n1602;
  assign n1604 = n1603 ^ n1498;
  assign n1634 = n1633 ^ n1604;
  assign n1594 = ~n721 & n821;
  assign n1595 = x73 & n824;
  assign n1596 = x72 & n898;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = x74 & n901;
  assign n1599 = n1597 & ~n1598;
  assign n1600 = ~n1594 & n1599;
  assign n1601 = n1600 ^ x14;
  assign n1635 = n1634 ^ n1601;
  assign n1591 = n1527 ^ n1487;
  assign n1592 = n1528 & n1591;
  assign n1593 = n1592 ^ n1487;
  assign n1636 = n1635 ^ n1593;
  assign n1583 = n596 & n956;
  assign n1584 = x75 & n673;
  assign n1585 = x76 & n601;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = x77 & n676;
  assign n1588 = n1586 & ~n1587;
  assign n1589 = ~n1583 & n1588;
  assign n1590 = n1589 ^ x11;
  assign n1637 = n1636 ^ n1590;
  assign n1580 = n1529 ^ n1476;
  assign n1581 = ~n1530 & ~n1580;
  assign n1582 = n1581 ^ n1476;
  assign n1638 = n1637 ^ n1582;
  assign n1572 = n399 & n1242;
  assign n1573 = x79 & n402;
  assign n1574 = x78 & n478;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = x80 & n470;
  assign n1577 = n1575 & ~n1576;
  assign n1578 = ~n1572 & n1577;
  assign n1579 = n1578 ^ x8;
  assign n1639 = n1638 ^ n1579;
  assign n1569 = n1531 ^ n1465;
  assign n1570 = n1532 & n1569;
  assign n1571 = n1570 ^ n1465;
  assign n1640 = n1639 ^ n1571;
  assign n1560 = n1226 ^ x83;
  assign n1561 = n239 & n1560;
  assign n1562 = x81 & n249;
  assign n1563 = x83 & n280;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = x82 & n242;
  assign n1566 = n1564 & ~n1565;
  assign n1567 = ~n1561 & n1566;
  assign n1568 = n1567 ^ x5;
  assign n1641 = n1640 ^ n1568;
  assign n1557 = n1533 ^ n1453;
  assign n1558 = ~n1534 & n1557;
  assign n1559 = n1558 ^ n1453;
  assign n1642 = n1641 ^ n1559;
  assign n1549 = x85 ^ x84;
  assign n1550 = ~n1444 & n1549;
  assign n1551 = n169 & ~n1550;
  assign n1552 = n1551 ^ x1;
  assign n1553 = n1552 ^ x86;
  assign n1541 = x85 ^ x2;
  assign n1542 = n1541 ^ x85;
  assign n1543 = n1541 ^ x84;
  assign n1544 = n1543 ^ n1541;
  assign n1545 = n1542 & ~n1544;
  assign n1546 = n1545 ^ n1541;
  assign n1547 = ~x1 & n1546;
  assign n1548 = n1547 ^ n1541;
  assign n1554 = n1553 ^ n1548;
  assign n1555 = ~x0 & n1554;
  assign n1556 = n1555 ^ n1553;
  assign n1643 = n1642 ^ n1556;
  assign n1538 = n1535 ^ n1437;
  assign n1539 = n1536 & ~n1538;
  assign n1540 = n1539 ^ n1437;
  assign n1644 = n1643 ^ n1540;
  assign n1731 = ~x20 & ~x21;
  assign n1742 = ~x22 & x23;
  assign n1743 = n1731 & n1742;
  assign n1744 = x64 & n1743;
  assign n1745 = x23 ^ x22;
  assign n1746 = n1507 & n1745;
  assign n1747 = n142 & n1746;
  assign n1748 = n1731 ^ n1625;
  assign n1749 = x22 & n1748;
  assign n1750 = n1749 ^ n1625;
  assign n1751 = ~n1747 & ~n1750;
  assign n1752 = x65 & ~n1751;
  assign n1753 = n152 & n1745;
  assign n1754 = x66 & n1507;
  assign n1755 = ~n1753 & n1754;
  assign n1756 = ~n1752 & ~n1755;
  assign n1757 = n1756 ^ x23;
  assign n1758 = x22 & x64;
  assign n1759 = n1625 & n1758;
  assign n1760 = n1756 & n1759;
  assign n1761 = n1757 & n1760;
  assign n1762 = n1761 ^ n1757;
  assign n1763 = ~n1744 & ~n1762;
  assign n1732 = ~n233 & ~n1731;
  assign n1733 = n1732 ^ n1625;
  assign n1734 = x64 ^ x22;
  assign n1735 = n1734 ^ x22;
  assign n1736 = n1732 ^ x22;
  assign n1737 = ~n1735 & n1736;
  assign n1738 = n1737 ^ x22;
  assign n1739 = ~n1733 & ~n1738;
  assign n1740 = n1739 ^ n1625;
  assign n1741 = x23 & n1740;
  assign n1764 = n1763 ^ n1741;
  assign n1723 = n420 & n1404;
  assign n1724 = x67 & n1514;
  assign n1725 = x69 & n1517;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = x68 & n1408;
  assign n1728 = n1726 & ~n1727;
  assign n1729 = ~n1723 & n1728;
  assign n1730 = n1729 ^ x20;
  assign n1765 = n1764 ^ n1730;
  assign n1720 = n1631 ^ n1620;
  assign n1721 = n1629 & ~n1720;
  assign n1722 = n1721 ^ n1631;
  assign n1766 = n1765 ^ n1722;
  assign n1712 = n575 & n1098;
  assign n1713 = x70 & n1198;
  assign n1714 = x72 & n1201;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = x71 & n1102;
  assign n1717 = n1715 & ~n1716;
  assign n1718 = ~n1712 & n1717;
  assign n1719 = n1718 ^ x17;
  assign n1767 = n1766 ^ n1719;
  assign n1709 = n1632 ^ n1604;
  assign n1710 = ~n1633 & ~n1709;
  assign n1711 = n1710 ^ n1604;
  assign n1768 = n1767 ^ n1711;
  assign n1701 = n789 & n821;
  assign n1702 = x73 & n898;
  assign n1703 = x75 & n901;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = x74 & n824;
  assign n1706 = n1704 & ~n1705;
  assign n1707 = ~n1701 & n1706;
  assign n1708 = n1707 ^ x14;
  assign n1769 = n1768 ^ n1708;
  assign n1698 = n1634 ^ n1593;
  assign n1699 = n1635 & n1698;
  assign n1700 = n1699 ^ n1593;
  assign n1770 = n1769 ^ n1700;
  assign n1690 = n596 & n1041;
  assign n1691 = x76 & n673;
  assign n1692 = x77 & n601;
  assign n1693 = ~n1691 & ~n1692;
  assign n1694 = x78 & n676;
  assign n1695 = n1693 & ~n1694;
  assign n1696 = ~n1690 & n1695;
  assign n1697 = n1696 ^ x11;
  assign n1771 = n1770 ^ n1697;
  assign n1687 = n1636 ^ n1582;
  assign n1688 = ~n1637 & ~n1687;
  assign n1689 = n1688 ^ n1582;
  assign n1772 = n1771 ^ n1689;
  assign n1679 = n399 & n1340;
  assign n1680 = x79 & n478;
  assign n1681 = x81 & n470;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = x80 & n402;
  assign n1684 = n1682 & ~n1683;
  assign n1685 = ~n1679 & n1684;
  assign n1686 = n1685 ^ x8;
  assign n1773 = n1772 ^ n1686;
  assign n1676 = n1638 ^ n1571;
  assign n1677 = n1639 & n1676;
  assign n1678 = n1677 ^ n1571;
  assign n1774 = n1773 ^ n1678;
  assign n1667 = n1330 ^ x84;
  assign n1668 = n239 & n1667;
  assign n1669 = x82 & n249;
  assign n1670 = x84 & n280;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = x83 & n242;
  assign n1673 = n1671 & ~n1672;
  assign n1674 = ~n1668 & n1673;
  assign n1675 = n1674 ^ x5;
  assign n1775 = n1774 ^ n1675;
  assign n1664 = n1640 ^ n1559;
  assign n1665 = ~n1641 & n1664;
  assign n1666 = n1665 ^ n1559;
  assign n1776 = n1775 ^ n1666;
  assign n1653 = x86 ^ x2;
  assign n1654 = n1653 ^ x86;
  assign n1655 = n1653 ^ x85;
  assign n1656 = n1655 ^ n1653;
  assign n1657 = n1654 & ~n1656;
  assign n1658 = n1657 ^ n1653;
  assign n1659 = ~x1 & n1658;
  assign n1660 = n1659 ^ n1653;
  assign n1648 = x86 ^ x85;
  assign n1649 = ~n1550 & n1648;
  assign n1650 = n169 & ~n1649;
  assign n1651 = n1650 ^ x1;
  assign n1652 = n1651 ^ x87;
  assign n1661 = n1660 ^ n1652;
  assign n1662 = ~x0 & n1661;
  assign n1663 = n1662 ^ n1652;
  assign n1777 = n1776 ^ n1663;
  assign n1645 = n1642 ^ n1540;
  assign n1646 = n1643 & ~n1645;
  assign n1647 = n1646 ^ n1540;
  assign n1778 = n1777 ^ n1647;
  assign n1882 = n1741 & n1763;
  assign n1867 = n1625 ^ x23;
  assign n1868 = n1867 ^ n1625;
  assign n1869 = n1748 & n1868;
  assign n1870 = n1869 ^ n1625;
  assign n1871 = n1745 & n1870;
  assign n1872 = x65 & n1871;
  assign n1873 = n1507 & ~n1745;
  assign n1874 = x67 & n1873;
  assign n1875 = ~n1872 & ~n1874;
  assign n1876 = x66 & n1750;
  assign n1877 = n1875 & ~n1876;
  assign n1878 = n285 & n1746;
  assign n1879 = n1877 & ~n1878;
  assign n1880 = n1879 ^ x23;
  assign n1865 = x24 ^ x23;
  assign n1866 = x64 & n1865;
  assign n1881 = n1880 ^ n1866;
  assign n1883 = n1882 ^ n1881;
  assign n1857 = n458 & n1404;
  assign n1858 = x68 & n1514;
  assign n1859 = x69 & n1408;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = x70 & n1517;
  assign n1862 = n1860 & ~n1861;
  assign n1863 = ~n1857 & n1862;
  assign n1864 = n1863 ^ x20;
  assign n1884 = n1883 ^ n1864;
  assign n1854 = n1764 ^ n1722;
  assign n1855 = n1765 & n1854;
  assign n1856 = n1855 ^ n1722;
  assign n1885 = n1884 ^ n1856;
  assign n1846 = ~n653 & n1098;
  assign n1847 = x71 & n1198;
  assign n1848 = x73 & n1201;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = x72 & n1102;
  assign n1851 = n1849 & ~n1850;
  assign n1852 = ~n1846 & n1851;
  assign n1853 = n1852 ^ x17;
  assign n1886 = n1885 ^ n1853;
  assign n1843 = n1766 ^ n1711;
  assign n1844 = ~n1767 & ~n1843;
  assign n1845 = n1844 ^ n1711;
  assign n1887 = n1886 ^ n1845;
  assign n1835 = n821 & n870;
  assign n1836 = x74 & n898;
  assign n1837 = x75 & n824;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = x76 & n901;
  assign n1840 = n1838 & ~n1839;
  assign n1841 = ~n1835 & n1840;
  assign n1842 = n1841 ^ x14;
  assign n1888 = n1887 ^ n1842;
  assign n1832 = n1768 ^ n1700;
  assign n1833 = n1769 & n1832;
  assign n1834 = n1833 ^ n1700;
  assign n1889 = n1888 ^ n1834;
  assign n1824 = n596 & n1149;
  assign n1825 = x77 & n673;
  assign n1826 = x79 & n676;
  assign n1827 = ~n1825 & ~n1826;
  assign n1828 = x78 & n601;
  assign n1829 = n1827 & ~n1828;
  assign n1830 = ~n1824 & n1829;
  assign n1831 = n1830 ^ x11;
  assign n1890 = n1889 ^ n1831;
  assign n1821 = n1770 ^ n1689;
  assign n1822 = ~n1771 & ~n1821;
  assign n1823 = n1822 ^ n1689;
  assign n1891 = n1890 ^ n1823;
  assign n1813 = n399 & n1454;
  assign n1814 = x80 & n478;
  assign n1815 = x81 & n402;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = x82 & n470;
  assign n1818 = n1816 & ~n1817;
  assign n1819 = ~n1813 & n1818;
  assign n1820 = n1819 ^ x8;
  assign n1892 = n1891 ^ n1820;
  assign n1810 = n1772 ^ n1678;
  assign n1811 = n1773 & n1810;
  assign n1812 = n1811 ^ n1678;
  assign n1893 = n1892 ^ n1812;
  assign n1801 = n1444 ^ x85;
  assign n1802 = n239 & n1801;
  assign n1803 = x83 & n249;
  assign n1804 = x84 & n242;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = x85 & n280;
  assign n1807 = n1805 & ~n1806;
  assign n1808 = ~n1802 & n1807;
  assign n1809 = n1808 ^ x5;
  assign n1894 = n1893 ^ n1809;
  assign n1798 = n1774 ^ n1666;
  assign n1799 = ~n1775 & n1798;
  assign n1800 = n1799 ^ n1666;
  assign n1895 = n1894 ^ n1800;
  assign n1790 = x87 ^ x86;
  assign n1791 = ~n1649 & n1790;
  assign n1792 = n169 & ~n1791;
  assign n1793 = n1792 ^ x1;
  assign n1794 = n1793 ^ x88;
  assign n1782 = x87 ^ x2;
  assign n1783 = n1782 ^ x87;
  assign n1784 = n1782 ^ x86;
  assign n1785 = n1784 ^ n1782;
  assign n1786 = n1783 & ~n1785;
  assign n1787 = n1786 ^ n1782;
  assign n1788 = ~x1 & n1787;
  assign n1789 = n1788 ^ n1782;
  assign n1795 = n1794 ^ n1789;
  assign n1796 = ~x0 & n1795;
  assign n1797 = n1796 ^ n1794;
  assign n1896 = n1895 ^ n1797;
  assign n1779 = n1776 ^ n1647;
  assign n1780 = n1777 & ~n1779;
  assign n1781 = n1780 ^ n1647;
  assign n1897 = n1896 ^ n1781;
  assign n2001 = ~n1866 & ~n1882;
  assign n2002 = ~n1880 & ~n2001;
  assign n1992 = n321 & n1746;
  assign n1993 = x66 & n1871;
  assign n1994 = x68 & n1873;
  assign n1995 = ~n1993 & ~n1994;
  assign n1996 = x67 & n1750;
  assign n1997 = n1995 & ~n1996;
  assign n1998 = ~n1992 & n1997;
  assign n1999 = n1998 ^ x23;
  assign n1987 = x65 ^ x24;
  assign n1988 = n1865 & ~n1987;
  assign n1989 = n1988 ^ x23;
  assign n1990 = n1989 ^ x25;
  assign n1984 = x23 & x24;
  assign n1985 = n1984 ^ x25;
  assign n1986 = ~x64 & n1985;
  assign n1991 = n1990 ^ n1986;
  assign n2000 = n1999 ^ n1991;
  assign n2003 = n2002 ^ n2000;
  assign n1976 = n517 & n1404;
  assign n1977 = x69 & n1514;
  assign n1978 = x70 & n1408;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = x71 & n1517;
  assign n1981 = n1979 & ~n1980;
  assign n1982 = ~n1976 & n1981;
  assign n1983 = n1982 ^ x20;
  assign n2004 = n2003 ^ n1983;
  assign n1973 = n1883 ^ n1856;
  assign n1974 = ~n1884 & ~n1973;
  assign n1975 = n1974 ^ n1856;
  assign n2005 = n2004 ^ n1975;
  assign n1965 = ~n721 & n1098;
  assign n1966 = x73 & n1102;
  assign n1967 = x72 & n1198;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = x74 & n1201;
  assign n1970 = n1968 & ~n1969;
  assign n1971 = ~n1965 & n1970;
  assign n1972 = n1971 ^ x17;
  assign n2006 = n2005 ^ n1972;
  assign n1962 = n1885 ^ n1845;
  assign n1963 = n1886 & n1962;
  assign n1964 = n1963 ^ n1845;
  assign n2007 = n2006 ^ n1964;
  assign n1954 = n821 & n956;
  assign n1955 = x75 & n898;
  assign n1956 = x76 & n824;
  assign n1957 = ~n1955 & ~n1956;
  assign n1958 = x77 & n901;
  assign n1959 = n1957 & ~n1958;
  assign n1960 = ~n1954 & n1959;
  assign n1961 = n1960 ^ x14;
  assign n2008 = n2007 ^ n1961;
  assign n1951 = n1887 ^ n1834;
  assign n1952 = ~n1888 & ~n1951;
  assign n1953 = n1952 ^ n1834;
  assign n2009 = n2008 ^ n1953;
  assign n1943 = n596 & n1242;
  assign n1944 = x78 & n673;
  assign n1945 = x79 & n601;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = x80 & n676;
  assign n1948 = n1946 & ~n1947;
  assign n1949 = ~n1943 & n1948;
  assign n1950 = n1949 ^ x11;
  assign n2010 = n2009 ^ n1950;
  assign n1940 = n1889 ^ n1823;
  assign n1941 = n1890 & n1940;
  assign n1942 = n1941 ^ n1823;
  assign n2011 = n2010 ^ n1942;
  assign n1932 = n399 & n1560;
  assign n1933 = x81 & n478;
  assign n1934 = x82 & n402;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = x83 & n470;
  assign n1937 = n1935 & ~n1936;
  assign n1938 = ~n1932 & n1937;
  assign n1939 = n1938 ^ x8;
  assign n2012 = n2011 ^ n1939;
  assign n1929 = n1891 ^ n1812;
  assign n1930 = ~n1892 & ~n1929;
  assign n1931 = n1930 ^ n1812;
  assign n2013 = n2012 ^ n1931;
  assign n1920 = n1550 ^ x86;
  assign n1921 = n239 & n1920;
  assign n1922 = x84 & n249;
  assign n1923 = x86 & n280;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = x85 & n242;
  assign n1926 = n1924 & ~n1925;
  assign n1927 = ~n1921 & n1926;
  assign n1928 = n1927 ^ x5;
  assign n2014 = n2013 ^ n1928;
  assign n1917 = n1893 ^ n1800;
  assign n1918 = n1894 & ~n1917;
  assign n1919 = n1918 ^ n1800;
  assign n2015 = n2014 ^ n1919;
  assign n1909 = x88 ^ x87;
  assign n1910 = ~n1791 & n1909;
  assign n1911 = n169 & ~n1910;
  assign n1912 = n1911 ^ x1;
  assign n1913 = n1912 ^ x89;
  assign n1901 = x88 ^ x2;
  assign n1902 = n1901 ^ x88;
  assign n1903 = n1901 ^ x87;
  assign n1904 = n1903 ^ n1901;
  assign n1905 = n1902 & ~n1904;
  assign n1906 = n1905 ^ n1901;
  assign n1907 = ~x1 & n1906;
  assign n1908 = n1907 ^ n1901;
  assign n1914 = n1913 ^ n1908;
  assign n1915 = ~x0 & n1914;
  assign n1916 = n1915 ^ n1913;
  assign n2016 = n2015 ^ n1916;
  assign n1898 = n1895 ^ n1781;
  assign n1899 = ~n1896 & n1898;
  assign n1900 = n1899 ^ n1781;
  assign n2017 = n2016 ^ n1900;
  assign n2135 = n789 & n1098;
  assign n2136 = x74 & n1102;
  assign n2137 = x73 & n1198;
  assign n2138 = ~n2136 & ~n2137;
  assign n2139 = x75 & n1201;
  assign n2140 = n2138 & ~n2139;
  assign n2141 = ~n2135 & n2140;
  assign n2142 = n2141 ^ x17;
  assign n2132 = n2005 ^ n1964;
  assign n2133 = n2006 & n2132;
  assign n2134 = n2133 ^ n1964;
  assign n2143 = n2142 ^ n2134;
  assign n2120 = n420 & n1746;
  assign n2121 = x67 & n1871;
  assign n2122 = x69 & n1873;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = x68 & n1750;
  assign n2125 = n2123 & ~n2124;
  assign n2126 = ~n2120 & n2125;
  assign n2127 = n2126 ^ x23;
  assign n2101 = x26 ^ x25;
  assign n2102 = n1865 & n2101;
  assign n2103 = n142 & n2102;
  assign n2104 = x25 & ~n1865;
  assign n2105 = n2104 ^ n1984;
  assign n2106 = ~n2103 & ~n2105;
  assign n2107 = x65 & ~n2106;
  assign n2108 = n1984 ^ x26;
  assign n2109 = n2108 ^ n1984;
  assign n2110 = ~n1865 & n2109;
  assign n2111 = n2110 ^ n1984;
  assign n2112 = n2101 & n2111;
  assign n2113 = x64 & n2112;
  assign n2114 = n152 & n2101;
  assign n2115 = x66 & n1865;
  assign n2116 = ~n2114 & n2115;
  assign n2117 = ~n2113 & ~n2116;
  assign n2118 = ~n2107 & n2117;
  assign n2095 = x25 ^ x23;
  assign n2096 = x64 & n2095;
  assign n2097 = n2096 ^ n233;
  assign n2098 = ~n1865 & ~n2097;
  assign n2099 = n2098 ^ n233;
  assign n2100 = x26 & ~n2099;
  assign n2119 = n2118 ^ n2100;
  assign n2128 = n2127 ^ n2119;
  assign n2092 = n2002 ^ n1999;
  assign n2093 = n2000 & ~n2092;
  assign n2094 = n2093 ^ n2002;
  assign n2129 = n2128 ^ n2094;
  assign n2084 = n575 & n1404;
  assign n2085 = x70 & n1514;
  assign n2086 = x72 & n1517;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = x71 & n1408;
  assign n2089 = n2087 & ~n2088;
  assign n2090 = ~n2084 & n2089;
  assign n2091 = n2090 ^ x20;
  assign n2130 = n2129 ^ n2091;
  assign n2081 = n2003 ^ n1975;
  assign n2082 = ~n2004 & ~n2081;
  assign n2083 = n2082 ^ n1975;
  assign n2131 = n2130 ^ n2083;
  assign n2144 = n2143 ^ n2131;
  assign n2073 = n821 & n1041;
  assign n2074 = x76 & n898;
  assign n2075 = x77 & n824;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = x78 & n901;
  assign n2078 = n2076 & ~n2077;
  assign n2079 = ~n2073 & n2078;
  assign n2080 = n2079 ^ x14;
  assign n2145 = n2144 ^ n2080;
  assign n2070 = n2007 ^ n1953;
  assign n2071 = ~n2008 & ~n2070;
  assign n2072 = n2071 ^ n1953;
  assign n2146 = n2145 ^ n2072;
  assign n2062 = n596 & n1340;
  assign n2063 = x79 & n673;
  assign n2064 = x81 & n676;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = x80 & n601;
  assign n2067 = n2065 & ~n2066;
  assign n2068 = ~n2062 & n2067;
  assign n2069 = n2068 ^ x11;
  assign n2147 = n2146 ^ n2069;
  assign n2059 = n2009 ^ n1942;
  assign n2060 = n2010 & n2059;
  assign n2061 = n2060 ^ n1942;
  assign n2148 = n2147 ^ n2061;
  assign n2051 = n399 & n1667;
  assign n2052 = x82 & n478;
  assign n2053 = x84 & n470;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = x83 & n402;
  assign n2056 = n2054 & ~n2055;
  assign n2057 = ~n2051 & n2056;
  assign n2058 = n2057 ^ x8;
  assign n2149 = n2148 ^ n2058;
  assign n2048 = n2011 ^ n1931;
  assign n2049 = ~n2012 & ~n2048;
  assign n2050 = n2049 ^ n1931;
  assign n2150 = n2149 ^ n2050;
  assign n2039 = n1649 ^ x87;
  assign n2040 = n239 & n2039;
  assign n2041 = x85 & n249;
  assign n2042 = x87 & n280;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = x86 & n242;
  assign n2045 = n2043 & ~n2044;
  assign n2046 = ~n2040 & n2045;
  assign n2047 = n2046 ^ x5;
  assign n2151 = n2150 ^ n2047;
  assign n2036 = n2013 ^ n1919;
  assign n2037 = n2014 & ~n2036;
  assign n2038 = n2037 ^ n1919;
  assign n2152 = n2151 ^ n2038;
  assign n2028 = x89 ^ x88;
  assign n2029 = ~n1910 & n2028;
  assign n2030 = n169 & ~n2029;
  assign n2031 = n2030 ^ x1;
  assign n2032 = n2031 ^ x90;
  assign n2021 = x2 & ~x88;
  assign n2022 = n2021 ^ x1;
  assign n2023 = n2022 ^ n2021;
  assign n2024 = x89 ^ x2;
  assign n2025 = n2024 ^ n2021;
  assign n2026 = n2023 & n2025;
  assign n2027 = n2026 ^ n2021;
  assign n2033 = n2032 ^ n2027;
  assign n2034 = ~x0 & n2033;
  assign n2035 = n2034 ^ n2032;
  assign n2153 = n2152 ^ n2035;
  assign n2018 = n2015 ^ n1900;
  assign n2019 = ~n2016 & n2018;
  assign n2020 = n2019 ^ n1900;
  assign n2154 = n2153 ^ n2020;
  assign n2260 = n458 & n1746;
  assign n2261 = x68 & n1871;
  assign n2262 = x70 & n1873;
  assign n2263 = ~n2261 & ~n2262;
  assign n2264 = x69 & n1750;
  assign n2265 = n2263 & ~n2264;
  assign n2266 = ~n2260 & n2265;
  assign n2267 = n2266 ^ x23;
  assign n2256 = x26 & n2099;
  assign n2257 = n2118 & n2256;
  assign n2254 = x27 ^ x26;
  assign n2255 = x64 & n2254;
  assign n2258 = n2257 ^ n2255;
  assign n2243 = x65 & n2112;
  assign n2244 = x66 & n2105;
  assign n2245 = ~n2243 & ~n2244;
  assign n2246 = n285 ^ x67;
  assign n2247 = n2101 ^ n285;
  assign n2248 = n2247 ^ n285;
  assign n2249 = n2246 & ~n2248;
  assign n2250 = n2249 ^ n285;
  assign n2251 = n1865 & n2250;
  assign n2252 = n2245 & ~n2251;
  assign n2253 = n2252 ^ x26;
  assign n2259 = n2258 ^ n2253;
  assign n2268 = n2267 ^ n2259;
  assign n2240 = n2127 ^ n2094;
  assign n2241 = ~n2128 & ~n2240;
  assign n2242 = n2241 ^ n2094;
  assign n2269 = n2268 ^ n2242;
  assign n2232 = ~n653 & n1404;
  assign n2233 = x71 & n1514;
  assign n2234 = x73 & n1517;
  assign n2235 = ~n2233 & ~n2234;
  assign n2236 = x72 & n1408;
  assign n2237 = n2235 & ~n2236;
  assign n2238 = ~n2232 & n2237;
  assign n2239 = n2238 ^ x20;
  assign n2270 = n2269 ^ n2239;
  assign n2229 = n2129 ^ n2083;
  assign n2230 = n2130 & n2229;
  assign n2231 = n2230 ^ n2083;
  assign n2271 = n2270 ^ n2231;
  assign n2221 = n870 & n1098;
  assign n2222 = x74 & n1198;
  assign n2223 = x76 & n1201;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = x75 & n1102;
  assign n2226 = n2224 & ~n2225;
  assign n2227 = ~n2221 & n2226;
  assign n2228 = n2227 ^ x17;
  assign n2272 = n2271 ^ n2228;
  assign n2218 = n2142 ^ n2131;
  assign n2219 = ~n2143 & ~n2218;
  assign n2220 = n2219 ^ n2134;
  assign n2273 = n2272 ^ n2220;
  assign n2210 = n821 & n1149;
  assign n2211 = x77 & n898;
  assign n2212 = x79 & n901;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = x78 & n824;
  assign n2215 = n2213 & ~n2214;
  assign n2216 = ~n2210 & n2215;
  assign n2217 = n2216 ^ x14;
  assign n2274 = n2273 ^ n2217;
  assign n2207 = n2144 ^ n2072;
  assign n2208 = n2145 & n2207;
  assign n2209 = n2208 ^ n2072;
  assign n2275 = n2274 ^ n2209;
  assign n2199 = n596 & n1454;
  assign n2200 = x80 & n673;
  assign n2201 = x81 & n601;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = x82 & n676;
  assign n2204 = n2202 & ~n2203;
  assign n2205 = ~n2199 & n2204;
  assign n2206 = n2205 ^ x11;
  assign n2276 = n2275 ^ n2206;
  assign n2196 = n2146 ^ n2061;
  assign n2197 = ~n2147 & ~n2196;
  assign n2198 = n2197 ^ n2061;
  assign n2277 = n2276 ^ n2198;
  assign n2188 = n399 & n1801;
  assign n2189 = x83 & n478;
  assign n2190 = x84 & n402;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = x85 & n470;
  assign n2193 = n2191 & ~n2192;
  assign n2194 = ~n2188 & n2193;
  assign n2195 = n2194 ^ x8;
  assign n2278 = n2277 ^ n2195;
  assign n2185 = n2148 ^ n2050;
  assign n2186 = n2149 & n2185;
  assign n2187 = n2186 ^ n2050;
  assign n2279 = n2278 ^ n2187;
  assign n2176 = n1791 ^ x88;
  assign n2177 = n239 & n2176;
  assign n2178 = x86 & n249;
  assign n2179 = x87 & n242;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = x88 & n280;
  assign n2182 = n2180 & ~n2181;
  assign n2183 = ~n2177 & n2182;
  assign n2184 = n2183 ^ x5;
  assign n2280 = n2279 ^ n2184;
  assign n2173 = n2150 ^ n2038;
  assign n2174 = ~n2151 & n2173;
  assign n2175 = n2174 ^ n2038;
  assign n2281 = n2280 ^ n2175;
  assign n2165 = x90 ^ x89;
  assign n2166 = ~n2029 & n2165;
  assign n2167 = n169 & ~n2166;
  assign n2168 = n2167 ^ x1;
  assign n2169 = n2168 ^ x91;
  assign n2158 = x2 & ~x89;
  assign n2159 = n2158 ^ x1;
  assign n2160 = n2159 ^ n2158;
  assign n2161 = x90 ^ x2;
  assign n2162 = n2161 ^ n2158;
  assign n2163 = n2160 & n2162;
  assign n2164 = n2163 ^ n2158;
  assign n2170 = n2169 ^ n2164;
  assign n2171 = ~x0 & n2170;
  assign n2172 = n2171 ^ n2169;
  assign n2282 = n2281 ^ n2172;
  assign n2155 = n2152 ^ n2020;
  assign n2156 = n2153 & ~n2155;
  assign n2157 = n2156 ^ n2020;
  assign n2283 = n2282 ^ n2157;
  assign n2398 = n517 & n1746;
  assign n2399 = x70 & n1750;
  assign n2400 = x69 & n1871;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = x71 & n1873;
  assign n2403 = n2401 & ~n2402;
  assign n2404 = ~n2398 & n2403;
  assign n2405 = n2404 ^ x23;
  assign n2395 = ~n2255 & ~n2257;
  assign n2396 = ~n2253 & ~n2395;
  assign n2390 = x26 & x27;
  assign n2391 = n2390 ^ x28;
  assign n2392 = ~x64 & n2391;
  assign n2386 = x65 ^ x27;
  assign n2387 = n2254 & ~n2386;
  assign n2388 = n2387 ^ x26;
  assign n2389 = n2388 ^ x28;
  assign n2393 = n2392 ^ n2389;
  assign n2377 = n321 & n2102;
  assign n2378 = x66 & n2112;
  assign n2379 = x67 & n2105;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = n1865 & ~n2101;
  assign n2382 = x68 & n2381;
  assign n2383 = n2380 & ~n2382;
  assign n2384 = ~n2377 & n2383;
  assign n2385 = n2384 ^ x26;
  assign n2394 = n2393 ^ n2385;
  assign n2397 = n2396 ^ n2394;
  assign n2406 = n2405 ^ n2397;
  assign n2374 = n2267 ^ n2242;
  assign n2375 = ~n2268 & ~n2374;
  assign n2376 = n2375 ^ n2242;
  assign n2407 = n2406 ^ n2376;
  assign n2366 = ~n721 & n1404;
  assign n2367 = x73 & n1408;
  assign n2368 = x74 & n1517;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = x72 & n1514;
  assign n2371 = n2369 & ~n2370;
  assign n2372 = ~n2366 & n2371;
  assign n2373 = n2372 ^ x20;
  assign n2408 = n2407 ^ n2373;
  assign n2363 = n2269 ^ n2231;
  assign n2364 = n2270 & n2363;
  assign n2365 = n2364 ^ n2231;
  assign n2409 = n2408 ^ n2365;
  assign n2355 = n956 & n1098;
  assign n2356 = x75 & n1198;
  assign n2357 = x76 & n1102;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = x77 & n1201;
  assign n2360 = n2358 & ~n2359;
  assign n2361 = ~n2355 & n2360;
  assign n2362 = n2361 ^ x17;
  assign n2410 = n2409 ^ n2362;
  assign n2352 = n2271 ^ n2220;
  assign n2353 = ~n2272 & ~n2352;
  assign n2354 = n2353 ^ n2220;
  assign n2411 = n2410 ^ n2354;
  assign n2344 = n821 & n1242;
  assign n2345 = x78 & n898;
  assign n2346 = x80 & n901;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = x79 & n824;
  assign n2349 = n2347 & ~n2348;
  assign n2350 = ~n2344 & n2349;
  assign n2351 = n2350 ^ x14;
  assign n2412 = n2411 ^ n2351;
  assign n2341 = n2273 ^ n2209;
  assign n2342 = n2274 & n2341;
  assign n2343 = n2342 ^ n2209;
  assign n2413 = n2412 ^ n2343;
  assign n2333 = n596 & n1560;
  assign n2334 = x81 & n673;
  assign n2335 = x82 & n601;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = x83 & n676;
  assign n2338 = n2336 & ~n2337;
  assign n2339 = ~n2333 & n2338;
  assign n2340 = n2339 ^ x11;
  assign n2414 = n2413 ^ n2340;
  assign n2330 = n2275 ^ n2198;
  assign n2331 = ~n2276 & ~n2330;
  assign n2332 = n2331 ^ n2198;
  assign n2415 = n2414 ^ n2332;
  assign n2322 = n399 & n1920;
  assign n2323 = x84 & n478;
  assign n2324 = x86 & n470;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = x85 & n402;
  assign n2327 = n2325 & ~n2326;
  assign n2328 = ~n2322 & n2327;
  assign n2329 = n2328 ^ x8;
  assign n2416 = n2415 ^ n2329;
  assign n2319 = n2277 ^ n2187;
  assign n2320 = n2278 & n2319;
  assign n2321 = n2320 ^ n2187;
  assign n2417 = n2416 ^ n2321;
  assign n2310 = n1910 ^ x89;
  assign n2311 = n239 & n2310;
  assign n2312 = x87 & n249;
  assign n2313 = x88 & n242;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = x89 & n280;
  assign n2316 = n2314 & ~n2315;
  assign n2317 = ~n2311 & n2316;
  assign n2318 = n2317 ^ x5;
  assign n2418 = n2417 ^ n2318;
  assign n2307 = n2279 ^ n2175;
  assign n2308 = ~n2280 & n2307;
  assign n2309 = n2308 ^ n2175;
  assign n2419 = n2418 ^ n2309;
  assign n2299 = x91 ^ x90;
  assign n2300 = ~n2166 & n2299;
  assign n2301 = n169 & ~n2300;
  assign n2302 = n2301 ^ x1;
  assign n2303 = n2302 ^ x92;
  assign n2287 = x91 ^ x2;
  assign n2288 = n2287 ^ x1;
  assign n2289 = n2288 ^ n2287;
  assign n2290 = n2289 ^ x0;
  assign n2291 = n2287 ^ x91;
  assign n2292 = n2291 ^ x90;
  assign n2293 = ~x90 & ~n2292;
  assign n2294 = n2293 ^ n2287;
  assign n2295 = n2294 ^ x90;
  assign n2296 = n2290 & ~n2295;
  assign n2297 = n2296 ^ n2293;
  assign n2298 = n2297 ^ x90;
  assign n2304 = n2303 ^ n2298;
  assign n2305 = ~x0 & ~n2304;
  assign n2306 = n2305 ^ n2303;
  assign n2420 = n2419 ^ n2306;
  assign n2284 = n2281 ^ n2157;
  assign n2285 = n2282 & ~n2284;
  assign n2286 = n2285 ^ n2157;
  assign n2421 = n2420 ^ n2286;
  assign n2558 = n575 & n1746;
  assign n2559 = x70 & n1871;
  assign n2560 = x72 & n1873;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = x71 & n1750;
  assign n2563 = n2561 & ~n2562;
  assign n2564 = ~n2558 & n2563;
  assign n2565 = n2564 ^ x23;
  assign n2526 = x29 ^ x28;
  assign n2527 = n2254 & n2526;
  assign n2528 = n142 & n2527;
  assign n2529 = x28 & ~n2254;
  assign n2530 = n2529 ^ n2390;
  assign n2531 = ~n2528 & ~n2530;
  assign n2532 = x65 & ~n2531;
  assign n2533 = n152 & n2526;
  assign n2534 = x66 & n2254;
  assign n2535 = ~n2533 & n2534;
  assign n2536 = ~n2532 & ~n2535;
  assign n2537 = ~x28 & x64;
  assign n2538 = x29 & ~n2537;
  assign n2539 = x28 ^ x26;
  assign n2540 = x64 & n2539;
  assign n2541 = n2540 ^ n233;
  assign n2542 = ~n2254 & ~n2541;
  assign n2543 = n2542 ^ n233;
  assign n2544 = n2538 & n2543;
  assign n2545 = n2536 & n2544;
  assign n2546 = n2536 ^ x29;
  assign n2547 = n2543 ^ n2536;
  assign n2548 = n2547 ^ n2543;
  assign n2549 = x28 & x64;
  assign n2550 = n2390 & n2549;
  assign n2551 = n2550 ^ n2543;
  assign n2552 = n2548 & n2551;
  assign n2553 = n2552 ^ n2543;
  assign n2554 = n2546 & ~n2553;
  assign n2555 = ~n2545 & ~n2554;
  assign n2518 = n420 & n2102;
  assign n2519 = x68 & n2105;
  assign n2520 = x67 & n2112;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = x69 & n2381;
  assign n2523 = n2521 & ~n2522;
  assign n2524 = ~n2518 & n2523;
  assign n2525 = n2524 ^ x26;
  assign n2556 = n2555 ^ n2525;
  assign n2515 = n2396 ^ n2385;
  assign n2516 = n2394 & ~n2515;
  assign n2517 = n2516 ^ n2396;
  assign n2557 = n2556 ^ n2517;
  assign n2566 = n2565 ^ n2557;
  assign n2512 = n2405 ^ n2376;
  assign n2513 = ~n2406 & ~n2512;
  assign n2514 = n2513 ^ n2376;
  assign n2567 = n2566 ^ n2514;
  assign n2504 = n789 & n1404;
  assign n2505 = x74 & n1408;
  assign n2506 = x75 & n1517;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = x73 & n1514;
  assign n2509 = n2507 & ~n2508;
  assign n2510 = ~n2504 & n2509;
  assign n2511 = n2510 ^ x20;
  assign n2568 = n2567 ^ n2511;
  assign n2501 = n2407 ^ n2365;
  assign n2502 = n2408 & n2501;
  assign n2503 = n2502 ^ n2365;
  assign n2569 = n2568 ^ n2503;
  assign n2493 = n1041 & n1098;
  assign n2494 = x76 & n1198;
  assign n2495 = x77 & n1102;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = x78 & n1201;
  assign n2498 = n2496 & ~n2497;
  assign n2499 = ~n2493 & n2498;
  assign n2500 = n2499 ^ x17;
  assign n2570 = n2569 ^ n2500;
  assign n2490 = n2409 ^ n2354;
  assign n2491 = ~n2410 & ~n2490;
  assign n2492 = n2491 ^ n2354;
  assign n2571 = n2570 ^ n2492;
  assign n2482 = n821 & n1340;
  assign n2483 = x79 & n898;
  assign n2484 = x81 & n901;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = x80 & n824;
  assign n2487 = n2485 & ~n2486;
  assign n2488 = ~n2482 & n2487;
  assign n2489 = n2488 ^ x14;
  assign n2572 = n2571 ^ n2489;
  assign n2479 = n2411 ^ n2343;
  assign n2480 = n2412 & n2479;
  assign n2481 = n2480 ^ n2343;
  assign n2573 = n2572 ^ n2481;
  assign n2471 = n596 & n1667;
  assign n2472 = x82 & n673;
  assign n2473 = x83 & n601;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = x84 & n676;
  assign n2476 = n2474 & ~n2475;
  assign n2477 = ~n2471 & n2476;
  assign n2478 = n2477 ^ x11;
  assign n2574 = n2573 ^ n2478;
  assign n2468 = n2413 ^ n2332;
  assign n2469 = ~n2414 & ~n2468;
  assign n2470 = n2469 ^ n2332;
  assign n2575 = n2574 ^ n2470;
  assign n2460 = n399 & n2039;
  assign n2461 = x85 & n478;
  assign n2462 = x86 & n402;
  assign n2463 = ~n2461 & ~n2462;
  assign n2464 = x87 & n470;
  assign n2465 = n2463 & ~n2464;
  assign n2466 = ~n2460 & n2465;
  assign n2467 = n2466 ^ x8;
  assign n2576 = n2575 ^ n2467;
  assign n2457 = n2415 ^ n2321;
  assign n2458 = n2416 & n2457;
  assign n2459 = n2458 ^ n2321;
  assign n2577 = n2576 ^ n2459;
  assign n2448 = n2029 ^ x90;
  assign n2449 = n239 & n2448;
  assign n2450 = x88 & n249;
  assign n2451 = x89 & n242;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = x90 & n280;
  assign n2454 = n2452 & ~n2453;
  assign n2455 = ~n2449 & n2454;
  assign n2456 = n2455 ^ x5;
  assign n2578 = n2577 ^ n2456;
  assign n2445 = n2417 ^ n2309;
  assign n2446 = ~n2418 & n2445;
  assign n2447 = n2446 ^ n2309;
  assign n2579 = n2578 ^ n2447;
  assign n2437 = x92 ^ x91;
  assign n2438 = ~n2300 & n2437;
  assign n2439 = n169 & ~n2438;
  assign n2440 = n2439 ^ x1;
  assign n2441 = n2440 ^ x93;
  assign n2425 = x92 ^ x2;
  assign n2426 = n2425 ^ x1;
  assign n2427 = n2426 ^ n2425;
  assign n2428 = n2427 ^ x0;
  assign n2429 = n2425 ^ x92;
  assign n2430 = n2429 ^ x91;
  assign n2431 = ~x91 & ~n2430;
  assign n2432 = n2431 ^ n2425;
  assign n2433 = n2432 ^ x91;
  assign n2434 = n2428 & ~n2433;
  assign n2435 = n2434 ^ n2431;
  assign n2436 = n2435 ^ x91;
  assign n2442 = n2441 ^ n2436;
  assign n2443 = ~x0 & ~n2442;
  assign n2444 = n2443 ^ n2441;
  assign n2580 = n2579 ^ n2444;
  assign n2422 = n2419 ^ n2286;
  assign n2423 = n2420 & ~n2422;
  assign n2424 = n2423 ^ n2286;
  assign n2581 = n2580 ^ n2424;
  assign n2703 = n458 & n2102;
  assign n2704 = x68 & n2112;
  assign n2705 = x69 & n2105;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = x70 & n2381;
  assign n2708 = n2706 & ~n2707;
  assign n2709 = ~n2703 & n2708;
  assign n2710 = n2709 ^ x26;
  assign n2699 = x30 ^ x29;
  assign n2700 = x64 & n2699;
  assign n2701 = n2700 ^ n2545;
  assign n2685 = x66 & n2530;
  assign n2686 = n2390 ^ x29;
  assign n2687 = n2686 ^ n2390;
  assign n2688 = ~n2254 & n2687;
  assign n2689 = n2688 ^ n2390;
  assign n2690 = n2526 & n2689;
  assign n2691 = x65 & n2690;
  assign n2692 = ~n2685 & ~n2691;
  assign n2693 = n2254 & ~n2526;
  assign n2694 = x67 & n2693;
  assign n2695 = n2692 & ~n2694;
  assign n2696 = n285 & n2527;
  assign n2697 = n2695 & ~n2696;
  assign n2698 = n2697 ^ x29;
  assign n2702 = n2701 ^ n2698;
  assign n2711 = n2710 ^ n2702;
  assign n2682 = n2555 ^ n2517;
  assign n2683 = n2556 & n2682;
  assign n2684 = n2683 ^ n2517;
  assign n2712 = n2711 ^ n2684;
  assign n2674 = ~n653 & n1746;
  assign n2675 = x71 & n1871;
  assign n2676 = x73 & n1873;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = x72 & n1750;
  assign n2679 = n2677 & ~n2678;
  assign n2680 = ~n2674 & n2679;
  assign n2681 = n2680 ^ x23;
  assign n2713 = n2712 ^ n2681;
  assign n2671 = n2565 ^ n2514;
  assign n2672 = ~n2566 & ~n2671;
  assign n2673 = n2672 ^ n2514;
  assign n2714 = n2713 ^ n2673;
  assign n2663 = n870 & n1404;
  assign n2664 = x75 & n1408;
  assign n2665 = x74 & n1514;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = x76 & n1517;
  assign n2668 = n2666 & ~n2667;
  assign n2669 = ~n2663 & n2668;
  assign n2670 = n2669 ^ x20;
  assign n2715 = n2714 ^ n2670;
  assign n2660 = n2567 ^ n2503;
  assign n2661 = n2568 & n2660;
  assign n2662 = n2661 ^ n2503;
  assign n2716 = n2715 ^ n2662;
  assign n2652 = n1098 & n1149;
  assign n2653 = x77 & n1198;
  assign n2654 = x78 & n1102;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = x79 & n1201;
  assign n2657 = n2655 & ~n2656;
  assign n2658 = ~n2652 & n2657;
  assign n2659 = n2658 ^ x17;
  assign n2717 = n2716 ^ n2659;
  assign n2649 = n2569 ^ n2492;
  assign n2650 = ~n2570 & ~n2649;
  assign n2651 = n2650 ^ n2492;
  assign n2718 = n2717 ^ n2651;
  assign n2641 = n821 & n1454;
  assign n2642 = x80 & n898;
  assign n2643 = x81 & n824;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = x82 & n901;
  assign n2646 = n2644 & ~n2645;
  assign n2647 = ~n2641 & n2646;
  assign n2648 = n2647 ^ x14;
  assign n2719 = n2718 ^ n2648;
  assign n2638 = n2571 ^ n2481;
  assign n2639 = n2572 & n2638;
  assign n2640 = n2639 ^ n2481;
  assign n2720 = n2719 ^ n2640;
  assign n2630 = n596 & n1801;
  assign n2631 = x83 & n673;
  assign n2632 = x85 & n676;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = x84 & n601;
  assign n2635 = n2633 & ~n2634;
  assign n2636 = ~n2630 & n2635;
  assign n2637 = n2636 ^ x11;
  assign n2721 = n2720 ^ n2637;
  assign n2627 = n2573 ^ n2470;
  assign n2628 = ~n2574 & ~n2627;
  assign n2629 = n2628 ^ n2470;
  assign n2722 = n2721 ^ n2629;
  assign n2619 = n399 & n2176;
  assign n2620 = x86 & n478;
  assign n2621 = x87 & n402;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = x88 & n470;
  assign n2624 = n2622 & ~n2623;
  assign n2625 = ~n2619 & n2624;
  assign n2626 = n2625 ^ x8;
  assign n2723 = n2722 ^ n2626;
  assign n2616 = n2575 ^ n2459;
  assign n2617 = n2576 & n2616;
  assign n2618 = n2617 ^ n2459;
  assign n2724 = n2723 ^ n2618;
  assign n2607 = n2166 ^ x91;
  assign n2608 = n239 & n2607;
  assign n2609 = x89 & n249;
  assign n2610 = x91 & n280;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = x90 & n242;
  assign n2613 = n2611 & ~n2612;
  assign n2614 = ~n2608 & n2613;
  assign n2615 = n2614 ^ x5;
  assign n2725 = n2724 ^ n2615;
  assign n2604 = n2577 ^ n2447;
  assign n2605 = ~n2578 & n2604;
  assign n2606 = n2605 ^ n2447;
  assign n2726 = n2725 ^ n2606;
  assign n2593 = x93 ^ x2;
  assign n2594 = n2593 ^ x93;
  assign n2595 = n2593 ^ x92;
  assign n2596 = n2595 ^ n2593;
  assign n2597 = n2594 & ~n2596;
  assign n2598 = n2597 ^ n2593;
  assign n2599 = ~x1 & n2598;
  assign n2600 = n2599 ^ n2593;
  assign n2585 = x93 ^ x92;
  assign n2586 = x93 ^ x91;
  assign n2587 = ~n2300 & ~n2586;
  assign n2588 = n2585 & n2587;
  assign n2589 = n2588 ^ n2585;
  assign n2590 = n169 & ~n2589;
  assign n2591 = n2590 ^ x1;
  assign n2592 = n2591 ^ x94;
  assign n2601 = n2600 ^ n2592;
  assign n2602 = ~x0 & n2601;
  assign n2603 = n2602 ^ n2592;
  assign n2727 = n2726 ^ n2603;
  assign n2582 = n2579 ^ n2424;
  assign n2583 = n2580 & ~n2582;
  assign n2584 = n2583 ^ n2424;
  assign n2728 = n2727 ^ n2584;
  assign n2853 = n517 & n2102;
  assign n2854 = x70 & n2105;
  assign n2855 = x69 & n2112;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = x71 & n2381;
  assign n2858 = n2856 & ~n2857;
  assign n2859 = ~n2853 & n2858;
  assign n2860 = n2859 ^ x26;
  assign n2850 = n2710 ^ n2684;
  assign n2851 = ~n2711 & ~n2850;
  assign n2852 = n2851 ^ n2684;
  assign n2861 = n2860 ^ n2852;
  assign n2847 = ~n2545 & ~n2700;
  assign n2848 = ~n2698 & ~n2847;
  assign n2838 = n321 & n2527;
  assign n2839 = x66 & n2690;
  assign n2840 = x68 & n2693;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = x67 & n2530;
  assign n2843 = n2841 & ~n2842;
  assign n2844 = ~n2838 & n2843;
  assign n2845 = n2844 ^ x29;
  assign n2833 = x65 ^ x30;
  assign n2834 = n2699 & ~n2833;
  assign n2835 = n2834 ^ x29;
  assign n2836 = n2835 ^ x31;
  assign n2830 = x29 & x30;
  assign n2831 = n2830 ^ x31;
  assign n2832 = ~x64 & n2831;
  assign n2837 = n2836 ^ n2832;
  assign n2846 = n2845 ^ n2837;
  assign n2849 = n2848 ^ n2846;
  assign n2862 = n2861 ^ n2849;
  assign n2822 = ~n721 & n1746;
  assign n2823 = x73 & n1750;
  assign n2824 = x72 & n1871;
  assign n2825 = ~n2823 & ~n2824;
  assign n2826 = x74 & n1873;
  assign n2827 = n2825 & ~n2826;
  assign n2828 = ~n2822 & n2827;
  assign n2829 = n2828 ^ x23;
  assign n2863 = n2862 ^ n2829;
  assign n2819 = n2712 ^ n2673;
  assign n2820 = n2713 & n2819;
  assign n2821 = n2820 ^ n2673;
  assign n2864 = n2863 ^ n2821;
  assign n2811 = n956 & n1404;
  assign n2812 = x75 & n1514;
  assign n2813 = x76 & n1408;
  assign n2814 = ~n2812 & ~n2813;
  assign n2815 = x77 & n1517;
  assign n2816 = n2814 & ~n2815;
  assign n2817 = ~n2811 & n2816;
  assign n2818 = n2817 ^ x20;
  assign n2865 = n2864 ^ n2818;
  assign n2808 = n2714 ^ n2662;
  assign n2809 = ~n2715 & ~n2808;
  assign n2810 = n2809 ^ n2662;
  assign n2866 = n2865 ^ n2810;
  assign n2800 = n1098 & n1242;
  assign n2801 = x78 & n1198;
  assign n2802 = x79 & n1102;
  assign n2803 = ~n2801 & ~n2802;
  assign n2804 = x80 & n1201;
  assign n2805 = n2803 & ~n2804;
  assign n2806 = ~n2800 & n2805;
  assign n2807 = n2806 ^ x17;
  assign n2867 = n2866 ^ n2807;
  assign n2797 = n2716 ^ n2651;
  assign n2798 = n2717 & n2797;
  assign n2799 = n2798 ^ n2651;
  assign n2868 = n2867 ^ n2799;
  assign n2789 = n821 & n1560;
  assign n2790 = x81 & n898;
  assign n2791 = x82 & n824;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = x83 & n901;
  assign n2794 = n2792 & ~n2793;
  assign n2795 = ~n2789 & n2794;
  assign n2796 = n2795 ^ x14;
  assign n2869 = n2868 ^ n2796;
  assign n2786 = n2718 ^ n2640;
  assign n2787 = ~n2719 & ~n2786;
  assign n2788 = n2787 ^ n2640;
  assign n2870 = n2869 ^ n2788;
  assign n2778 = n596 & n1920;
  assign n2779 = x84 & n673;
  assign n2780 = x85 & n601;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = x86 & n676;
  assign n2783 = n2781 & ~n2782;
  assign n2784 = ~n2778 & n2783;
  assign n2785 = n2784 ^ x11;
  assign n2871 = n2870 ^ n2785;
  assign n2775 = n2720 ^ n2629;
  assign n2776 = n2721 & n2775;
  assign n2777 = n2776 ^ n2629;
  assign n2872 = n2871 ^ n2777;
  assign n2767 = n399 & n2310;
  assign n2768 = x87 & n478;
  assign n2769 = x88 & n402;
  assign n2770 = ~n2768 & ~n2769;
  assign n2771 = x89 & n470;
  assign n2772 = n2770 & ~n2771;
  assign n2773 = ~n2767 & n2772;
  assign n2774 = n2773 ^ x8;
  assign n2873 = n2872 ^ n2774;
  assign n2764 = n2722 ^ n2618;
  assign n2765 = ~n2723 & ~n2764;
  assign n2766 = n2765 ^ n2618;
  assign n2874 = n2873 ^ n2766;
  assign n2755 = n2300 ^ x92;
  assign n2756 = n239 & n2755;
  assign n2757 = x90 & n249;
  assign n2758 = x91 & n242;
  assign n2759 = ~n2757 & ~n2758;
  assign n2760 = x92 & n280;
  assign n2761 = n2759 & ~n2760;
  assign n2762 = ~n2756 & n2761;
  assign n2763 = n2762 ^ x5;
  assign n2875 = n2874 ^ n2763;
  assign n2752 = n2724 ^ n2606;
  assign n2753 = n2725 & ~n2752;
  assign n2754 = n2753 ^ n2606;
  assign n2876 = n2875 ^ n2754;
  assign n2744 = x94 ^ x93;
  assign n2745 = ~n2589 & n2744;
  assign n2746 = n169 & ~n2745;
  assign n2747 = n2746 ^ x1;
  assign n2748 = n2747 ^ x95;
  assign n2732 = x94 ^ x2;
  assign n2733 = n2732 ^ x1;
  assign n2734 = n2733 ^ n2732;
  assign n2735 = n2734 ^ x0;
  assign n2736 = n2732 ^ x94;
  assign n2737 = n2736 ^ x93;
  assign n2738 = ~x93 & ~n2737;
  assign n2739 = n2738 ^ n2732;
  assign n2740 = n2739 ^ x93;
  assign n2741 = n2735 & ~n2740;
  assign n2742 = n2741 ^ n2738;
  assign n2743 = n2742 ^ x93;
  assign n2749 = n2748 ^ n2743;
  assign n2750 = ~x0 & ~n2749;
  assign n2751 = n2750 ^ n2748;
  assign n2877 = n2876 ^ n2751;
  assign n2729 = n2726 ^ n2584;
  assign n2730 = ~n2727 & n2729;
  assign n2731 = n2730 ^ n2584;
  assign n2878 = n2877 ^ n2731;
  assign n3004 = ~x29 & ~x30;
  assign n3005 = ~x31 & x32;
  assign n3006 = n3004 & n3005;
  assign n3007 = x64 & n3006;
  assign n3008 = x32 ^ x31;
  assign n3009 = n2699 & n3008;
  assign n3010 = n142 & n3009;
  assign n3011 = n3004 ^ n2830;
  assign n3012 = x31 & n3011;
  assign n3013 = n3012 ^ n2830;
  assign n3014 = ~n3010 & ~n3013;
  assign n3015 = x65 & ~n3014;
  assign n3016 = n152 & n3008;
  assign n3017 = x66 & n2699;
  assign n3018 = ~n3016 & n3017;
  assign n3019 = ~n3015 & ~n3018;
  assign n3020 = n3019 ^ x32;
  assign n3021 = x31 & x64;
  assign n3022 = n2830 & n3021;
  assign n3023 = n3019 & n3022;
  assign n3024 = n3020 & n3023;
  assign n3025 = n3024 ^ n3020;
  assign n3026 = ~n3007 & ~n3025;
  assign n2998 = x31 ^ x29;
  assign n2999 = x64 & n2998;
  assign n3000 = n2999 ^ n233;
  assign n3001 = ~n2699 & ~n3000;
  assign n3002 = n3001 ^ n233;
  assign n3003 = x32 & n3002;
  assign n3027 = n3026 ^ n3003;
  assign n2990 = n420 & n2527;
  assign n2991 = x67 & n2690;
  assign n2992 = x69 & n2693;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = x68 & n2530;
  assign n2995 = n2993 & ~n2994;
  assign n2996 = ~n2990 & n2995;
  assign n2997 = n2996 ^ x29;
  assign n3028 = n3027 ^ n2997;
  assign n2987 = n2848 ^ n2845;
  assign n2988 = n2846 & ~n2987;
  assign n2989 = n2988 ^ n2848;
  assign n3029 = n3028 ^ n2989;
  assign n2979 = n575 & n2102;
  assign n2980 = x71 & n2105;
  assign n2981 = x70 & n2112;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = x72 & n2381;
  assign n2984 = n2982 & ~n2983;
  assign n2985 = ~n2979 & n2984;
  assign n2986 = n2985 ^ x26;
  assign n3030 = n3029 ^ n2986;
  assign n2976 = n2860 ^ n2849;
  assign n2977 = ~n2861 & ~n2976;
  assign n2978 = n2977 ^ n2852;
  assign n3031 = n3030 ^ n2978;
  assign n2968 = n789 & n1746;
  assign n2969 = x73 & n1871;
  assign n2970 = x74 & n1750;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = x75 & n1873;
  assign n2973 = n2971 & ~n2972;
  assign n2974 = ~n2968 & n2973;
  assign n2975 = n2974 ^ x23;
  assign n3032 = n3031 ^ n2975;
  assign n2965 = n2862 ^ n2821;
  assign n2966 = n2863 & n2965;
  assign n2967 = n2966 ^ n2821;
  assign n3033 = n3032 ^ n2967;
  assign n2957 = n1041 & n1404;
  assign n2958 = x76 & n1514;
  assign n2959 = x77 & n1408;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = x78 & n1517;
  assign n2962 = n2960 & ~n2961;
  assign n2963 = ~n2957 & n2962;
  assign n2964 = n2963 ^ x20;
  assign n3034 = n3033 ^ n2964;
  assign n2954 = n2864 ^ n2810;
  assign n2955 = ~n2865 & ~n2954;
  assign n2956 = n2955 ^ n2810;
  assign n3035 = n3034 ^ n2956;
  assign n2946 = n1098 & n1340;
  assign n2947 = x79 & n1198;
  assign n2948 = x80 & n1102;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = x81 & n1201;
  assign n2951 = n2949 & ~n2950;
  assign n2952 = ~n2946 & n2951;
  assign n2953 = n2952 ^ x17;
  assign n3036 = n3035 ^ n2953;
  assign n2943 = n2866 ^ n2799;
  assign n2944 = n2867 & n2943;
  assign n2945 = n2944 ^ n2799;
  assign n3037 = n3036 ^ n2945;
  assign n2935 = n821 & n1667;
  assign n2936 = x82 & n898;
  assign n2937 = x84 & n901;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = x83 & n824;
  assign n2940 = n2938 & ~n2939;
  assign n2941 = ~n2935 & n2940;
  assign n2942 = n2941 ^ x14;
  assign n3038 = n3037 ^ n2942;
  assign n2932 = n2868 ^ n2788;
  assign n2933 = ~n2869 & ~n2932;
  assign n2934 = n2933 ^ n2788;
  assign n3039 = n3038 ^ n2934;
  assign n2924 = n596 & n2039;
  assign n2925 = x85 & n673;
  assign n2926 = x87 & n676;
  assign n2927 = ~n2925 & ~n2926;
  assign n2928 = x86 & n601;
  assign n2929 = n2927 & ~n2928;
  assign n2930 = ~n2924 & n2929;
  assign n2931 = n2930 ^ x11;
  assign n3040 = n3039 ^ n2931;
  assign n2921 = n2870 ^ n2777;
  assign n2922 = n2871 & n2921;
  assign n2923 = n2922 ^ n2777;
  assign n3041 = n3040 ^ n2923;
  assign n2913 = n399 & n2448;
  assign n2914 = x89 & n402;
  assign n2915 = x88 & n478;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = x90 & n470;
  assign n2918 = n2916 & ~n2917;
  assign n2919 = ~n2913 & n2918;
  assign n2920 = n2919 ^ x8;
  assign n3042 = n3041 ^ n2920;
  assign n2910 = n2872 ^ n2766;
  assign n2911 = ~n2873 & ~n2910;
  assign n2912 = n2911 ^ n2766;
  assign n3043 = n3042 ^ n2912;
  assign n2901 = n2438 ^ x93;
  assign n2902 = n239 & n2901;
  assign n2903 = x91 & n249;
  assign n2904 = x92 & n242;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = x93 & n280;
  assign n2907 = n2905 & ~n2906;
  assign n2908 = ~n2902 & n2907;
  assign n2909 = n2908 ^ x5;
  assign n3044 = n3043 ^ n2909;
  assign n2898 = n2874 ^ n2754;
  assign n2899 = n2875 & ~n2898;
  assign n2900 = n2899 ^ n2754;
  assign n3045 = n3044 ^ n2900;
  assign n2890 = x95 ^ x94;
  assign n2891 = ~n2745 & n2890;
  assign n2892 = n169 & ~n2891;
  assign n2893 = n2892 ^ x1;
  assign n2894 = n2893 ^ x96;
  assign n2882 = x95 ^ x2;
  assign n2883 = n2882 ^ x95;
  assign n2884 = n2882 ^ x94;
  assign n2885 = n2884 ^ n2882;
  assign n2886 = n2883 & ~n2885;
  assign n2887 = n2886 ^ n2882;
  assign n2888 = ~x1 & n2887;
  assign n2889 = n2888 ^ n2882;
  assign n2895 = n2894 ^ n2889;
  assign n2896 = ~x0 & n2895;
  assign n2897 = n2896 ^ n2894;
  assign n3046 = n3045 ^ n2897;
  assign n2879 = n2876 ^ n2731;
  assign n2880 = ~n2877 & n2879;
  assign n2881 = n2880 ^ n2731;
  assign n3047 = n3046 ^ n2881;
  assign n3192 = n3003 & n3026;
  assign n3177 = n2830 ^ x32;
  assign n3178 = n3177 ^ n2830;
  assign n3179 = n3011 & n3178;
  assign n3180 = n3179 ^ n2830;
  assign n3181 = n3008 & n3180;
  assign n3182 = x65 & n3181;
  assign n3183 = n2699 & ~n3008;
  assign n3184 = x67 & n3183;
  assign n3185 = ~n3182 & ~n3184;
  assign n3186 = x66 & n3013;
  assign n3187 = n3185 & ~n3186;
  assign n3188 = n285 & n3009;
  assign n3189 = n3187 & ~n3188;
  assign n3190 = n3189 ^ x32;
  assign n3175 = x33 ^ x32;
  assign n3176 = x64 & n3175;
  assign n3191 = n3190 ^ n3176;
  assign n3193 = n3192 ^ n3191;
  assign n3167 = n458 & n2527;
  assign n3168 = x69 & n2530;
  assign n3169 = x68 & n2690;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = x70 & n2693;
  assign n3172 = n3170 & ~n3171;
  assign n3173 = ~n3167 & n3172;
  assign n3174 = n3173 ^ x29;
  assign n3194 = n3193 ^ n3174;
  assign n3164 = n3027 ^ n2989;
  assign n3165 = n3028 & n3164;
  assign n3166 = n3165 ^ n2989;
  assign n3195 = n3194 ^ n3166;
  assign n3156 = ~n653 & n2102;
  assign n3157 = x72 & n2105;
  assign n3158 = x71 & n2112;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = x73 & n2381;
  assign n3161 = n3159 & ~n3160;
  assign n3162 = ~n3156 & n3161;
  assign n3163 = n3162 ^ x26;
  assign n3196 = n3195 ^ n3163;
  assign n3153 = n3029 ^ n2978;
  assign n3154 = ~n3030 & ~n3153;
  assign n3155 = n3154 ^ n2978;
  assign n3197 = n3196 ^ n3155;
  assign n3145 = n870 & n1746;
  assign n3146 = x74 & n1871;
  assign n3147 = x76 & n1873;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = x75 & n1750;
  assign n3150 = n3148 & ~n3149;
  assign n3151 = ~n3145 & n3150;
  assign n3152 = n3151 ^ x23;
  assign n3198 = n3197 ^ n3152;
  assign n3142 = n3031 ^ n2967;
  assign n3143 = n3032 & n3142;
  assign n3144 = n3143 ^ n2967;
  assign n3199 = n3198 ^ n3144;
  assign n3134 = n1149 & n1404;
  assign n3135 = x77 & n1514;
  assign n3136 = x78 & n1408;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = x79 & n1517;
  assign n3139 = n3137 & ~n3138;
  assign n3140 = ~n3134 & n3139;
  assign n3141 = n3140 ^ x20;
  assign n3200 = n3199 ^ n3141;
  assign n3131 = n3033 ^ n2956;
  assign n3132 = ~n3034 & ~n3131;
  assign n3133 = n3132 ^ n2956;
  assign n3201 = n3200 ^ n3133;
  assign n3123 = n1098 & n1454;
  assign n3124 = x80 & n1198;
  assign n3125 = x81 & n1102;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = x82 & n1201;
  assign n3128 = n3126 & ~n3127;
  assign n3129 = ~n3123 & n3128;
  assign n3130 = n3129 ^ x17;
  assign n3202 = n3201 ^ n3130;
  assign n3120 = n3035 ^ n2945;
  assign n3121 = n3036 & n3120;
  assign n3122 = n3121 ^ n2945;
  assign n3203 = n3202 ^ n3122;
  assign n3112 = n821 & n1801;
  assign n3113 = x83 & n898;
  assign n3114 = x85 & n901;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = x84 & n824;
  assign n3117 = n3115 & ~n3116;
  assign n3118 = ~n3112 & n3117;
  assign n3119 = n3118 ^ x14;
  assign n3204 = n3203 ^ n3119;
  assign n3109 = n3037 ^ n2934;
  assign n3110 = ~n3038 & ~n3109;
  assign n3111 = n3110 ^ n2934;
  assign n3205 = n3204 ^ n3111;
  assign n3101 = n596 & n2176;
  assign n3102 = x86 & n673;
  assign n3103 = x87 & n601;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = x88 & n676;
  assign n3106 = n3104 & ~n3105;
  assign n3107 = ~n3101 & n3106;
  assign n3108 = n3107 ^ x11;
  assign n3206 = n3205 ^ n3108;
  assign n3098 = n3039 ^ n2923;
  assign n3099 = n3040 & n3098;
  assign n3100 = n3099 ^ n2923;
  assign n3207 = n3206 ^ n3100;
  assign n3090 = n399 & n2607;
  assign n3091 = x89 & n478;
  assign n3092 = x91 & n470;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = x90 & n402;
  assign n3095 = n3093 & ~n3094;
  assign n3096 = ~n3090 & n3095;
  assign n3097 = n3096 ^ x8;
  assign n3208 = n3207 ^ n3097;
  assign n3087 = n3041 ^ n2912;
  assign n3088 = ~n3042 & ~n3087;
  assign n3089 = n3088 ^ n2912;
  assign n3209 = n3208 ^ n3089;
  assign n3078 = n2589 ^ x94;
  assign n3079 = n239 & n3078;
  assign n3080 = x92 & n249;
  assign n3081 = x94 & n280;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = x93 & n242;
  assign n3084 = n3082 & ~n3083;
  assign n3085 = ~n3079 & n3084;
  assign n3086 = n3085 ^ x5;
  assign n3210 = n3209 ^ n3086;
  assign n3075 = n3043 ^ n2900;
  assign n3076 = n3044 & ~n3075;
  assign n3077 = n3076 ^ n2900;
  assign n3211 = n3210 ^ n3077;
  assign n3059 = x96 ^ x95;
  assign n3060 = x96 ^ x94;
  assign n3061 = n2745 ^ x94;
  assign n3062 = n3061 ^ x94;
  assign n3063 = n3062 ^ x94;
  assign n3064 = n3063 ^ x94;
  assign n3065 = ~n3060 & n3064;
  assign n3066 = n3065 ^ x94;
  assign n3067 = n3066 ^ x96;
  assign n3068 = n3059 & n3067;
  assign n3069 = n169 & ~n3068;
  assign n3070 = n3069 ^ x1;
  assign n3071 = n3070 ^ x97;
  assign n3051 = x96 ^ x2;
  assign n3052 = n3051 ^ x95;
  assign n3053 = n3052 ^ n3051;
  assign n3054 = n3051 ^ x96;
  assign n3055 = ~n3053 & n3054;
  assign n3056 = n3055 ^ n3051;
  assign n3057 = ~x1 & n3056;
  assign n3058 = n3057 ^ n3051;
  assign n3072 = n3071 ^ n3058;
  assign n3073 = ~x0 & n3072;
  assign n3074 = n3073 ^ n3071;
  assign n3212 = n3211 ^ n3074;
  assign n3048 = n3045 ^ n2881;
  assign n3049 = ~n3046 & n3048;
  assign n3050 = n3049 ^ n2881;
  assign n3213 = n3212 ^ n3050;
  assign n3361 = ~n3176 & ~n3192;
  assign n3362 = ~n3190 & ~n3361;
  assign n3356 = x32 & x33;
  assign n3357 = n3356 ^ x34;
  assign n3358 = ~x64 & n3357;
  assign n3352 = x65 ^ x33;
  assign n3353 = n3175 & ~n3352;
  assign n3354 = n3353 ^ x32;
  assign n3355 = n3354 ^ x34;
  assign n3359 = n3358 ^ n3355;
  assign n3344 = n321 & n3009;
  assign n3345 = x67 & n3013;
  assign n3346 = x66 & n3181;
  assign n3347 = ~n3345 & ~n3346;
  assign n3348 = x68 & n3183;
  assign n3349 = n3347 & ~n3348;
  assign n3350 = ~n3344 & n3349;
  assign n3351 = n3350 ^ x32;
  assign n3360 = n3359 ^ n3351;
  assign n3363 = n3362 ^ n3360;
  assign n3336 = n517 & n2527;
  assign n3337 = x69 & n2690;
  assign n3338 = x71 & n2693;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = x70 & n2530;
  assign n3341 = n3339 & ~n3340;
  assign n3342 = ~n3336 & n3341;
  assign n3343 = n3342 ^ x29;
  assign n3364 = n3363 ^ n3343;
  assign n3333 = n3193 ^ n3166;
  assign n3334 = ~n3194 & ~n3333;
  assign n3335 = n3334 ^ n3166;
  assign n3365 = n3364 ^ n3335;
  assign n3325 = ~n721 & n2102;
  assign n3326 = x73 & n2105;
  assign n3327 = x72 & n2112;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = x74 & n2381;
  assign n3330 = n3328 & ~n3329;
  assign n3331 = ~n3325 & n3330;
  assign n3332 = n3331 ^ x26;
  assign n3366 = n3365 ^ n3332;
  assign n3322 = n3195 ^ n3155;
  assign n3323 = n3196 & n3322;
  assign n3324 = n3323 ^ n3155;
  assign n3367 = n3366 ^ n3324;
  assign n3314 = n956 & n1746;
  assign n3315 = x75 & n1871;
  assign n3316 = x76 & n1750;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = x77 & n1873;
  assign n3319 = n3317 & ~n3318;
  assign n3320 = ~n3314 & n3319;
  assign n3321 = n3320 ^ x23;
  assign n3368 = n3367 ^ n3321;
  assign n3311 = n3197 ^ n3144;
  assign n3312 = ~n3198 & ~n3311;
  assign n3313 = n3312 ^ n3144;
  assign n3369 = n3368 ^ n3313;
  assign n3303 = n1242 & n1404;
  assign n3304 = x78 & n1514;
  assign n3305 = x79 & n1408;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = x80 & n1517;
  assign n3308 = n3306 & ~n3307;
  assign n3309 = ~n3303 & n3308;
  assign n3310 = n3309 ^ x20;
  assign n3370 = n3369 ^ n3310;
  assign n3300 = n3199 ^ n3133;
  assign n3301 = n3200 & n3300;
  assign n3302 = n3301 ^ n3133;
  assign n3371 = n3370 ^ n3302;
  assign n3292 = n1098 & n1560;
  assign n3293 = x82 & n1102;
  assign n3294 = x81 & n1198;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = x83 & n1201;
  assign n3297 = n3295 & ~n3296;
  assign n3298 = ~n3292 & n3297;
  assign n3299 = n3298 ^ x17;
  assign n3372 = n3371 ^ n3299;
  assign n3289 = n3201 ^ n3122;
  assign n3290 = ~n3202 & ~n3289;
  assign n3291 = n3290 ^ n3122;
  assign n3373 = n3372 ^ n3291;
  assign n3281 = n821 & n1920;
  assign n3282 = x84 & n898;
  assign n3283 = x85 & n824;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = x86 & n901;
  assign n3286 = n3284 & ~n3285;
  assign n3287 = ~n3281 & n3286;
  assign n3288 = n3287 ^ x14;
  assign n3374 = n3373 ^ n3288;
  assign n3278 = n3203 ^ n3111;
  assign n3279 = n3204 & n3278;
  assign n3280 = n3279 ^ n3111;
  assign n3375 = n3374 ^ n3280;
  assign n3270 = n596 & n2310;
  assign n3271 = x87 & n673;
  assign n3272 = x89 & n676;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = x88 & n601;
  assign n3275 = n3273 & ~n3274;
  assign n3276 = ~n3270 & n3275;
  assign n3277 = n3276 ^ x11;
  assign n3376 = n3375 ^ n3277;
  assign n3267 = n3205 ^ n3100;
  assign n3268 = ~n3206 & ~n3267;
  assign n3269 = n3268 ^ n3100;
  assign n3377 = n3376 ^ n3269;
  assign n3259 = n399 & n2755;
  assign n3260 = x90 & n478;
  assign n3261 = x91 & n402;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = x92 & n470;
  assign n3264 = n3262 & ~n3263;
  assign n3265 = ~n3259 & n3264;
  assign n3266 = n3265 ^ x8;
  assign n3378 = n3377 ^ n3266;
  assign n3256 = n3207 ^ n3089;
  assign n3257 = n3208 & n3256;
  assign n3258 = n3257 ^ n3089;
  assign n3379 = n3378 ^ n3258;
  assign n3247 = n2745 ^ x95;
  assign n3248 = n239 & n3247;
  assign n3249 = x93 & n249;
  assign n3250 = x94 & n242;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = x95 & n280;
  assign n3253 = n3251 & ~n3252;
  assign n3254 = ~n3248 & n3253;
  assign n3255 = n3254 ^ x5;
  assign n3380 = n3379 ^ n3255;
  assign n3244 = n3209 ^ n3077;
  assign n3245 = ~n3210 & n3244;
  assign n3246 = n3245 ^ n3077;
  assign n3381 = n3380 ^ n3246;
  assign n3218 = x97 ^ x96;
  assign n3219 = x97 ^ x94;
  assign n3220 = n3219 ^ n2745;
  assign n3221 = n3219 ^ n3059;
  assign n3222 = n3219 & n3221;
  assign n3223 = n3222 ^ n3219;
  assign n3224 = ~n3220 & n3223;
  assign n3225 = n3224 ^ n3222;
  assign n3226 = n3225 ^ n3219;
  assign n3227 = n3226 ^ n3059;
  assign n3228 = n3218 & n3227;
  assign n3229 = n3228 ^ x96;
  assign n3230 = n3229 ^ x97;
  assign n3231 = n169 & ~n3230;
  assign n3232 = n3231 ^ x1;
  assign n3233 = n3232 ^ x98;
  assign n3217 = ~x96 & n197;
  assign n3234 = n3233 ^ n3217;
  assign n3235 = n3234 ^ n3233;
  assign n3236 = x97 ^ x2;
  assign n3237 = x1 & n3236;
  assign n3238 = n3237 ^ n3233;
  assign n3239 = n3238 ^ n3233;
  assign n3240 = ~n3235 & ~n3239;
  assign n3241 = n3240 ^ n3233;
  assign n3242 = ~x0 & ~n3241;
  assign n3243 = n3242 ^ n3233;
  assign n3382 = n3381 ^ n3243;
  assign n3214 = n3211 ^ n3050;
  assign n3215 = n3212 & ~n3214;
  assign n3216 = n3215 ^ n3050;
  assign n3383 = n3382 ^ n3216;
  assign n3517 = ~x32 & ~x33;
  assign n3518 = ~x34 & x35;
  assign n3519 = n3517 & n3518;
  assign n3520 = x64 & n3519;
  assign n3521 = x35 ^ x34;
  assign n3522 = n3175 & n3521;
  assign n3523 = n142 & n3522;
  assign n3524 = n3517 ^ n3356;
  assign n3525 = x34 & n3524;
  assign n3526 = n3525 ^ n3356;
  assign n3527 = ~n3523 & ~n3526;
  assign n3528 = x65 & ~n3527;
  assign n3529 = n152 & n3521;
  assign n3530 = x66 & n3175;
  assign n3531 = ~n3529 & n3530;
  assign n3532 = ~n3528 & ~n3531;
  assign n3533 = n3532 ^ x35;
  assign n3534 = x34 & x64;
  assign n3535 = n3356 & n3534;
  assign n3536 = n3532 & n3535;
  assign n3537 = n3533 & n3536;
  assign n3538 = n3537 ^ n3533;
  assign n3539 = ~n3520 & ~n3538;
  assign n3511 = x34 ^ x32;
  assign n3512 = x64 & n3511;
  assign n3513 = n3512 ^ n233;
  assign n3514 = ~n3175 & ~n3513;
  assign n3515 = n3514 ^ n233;
  assign n3516 = x35 & n3515;
  assign n3540 = n3539 ^ n3516;
  assign n3503 = n420 & n3009;
  assign n3504 = x68 & n3013;
  assign n3505 = x67 & n3181;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = x69 & n3183;
  assign n3508 = n3506 & ~n3507;
  assign n3509 = ~n3503 & n3508;
  assign n3510 = n3509 ^ x32;
  assign n3541 = n3540 ^ n3510;
  assign n3500 = n3362 ^ n3351;
  assign n3501 = n3360 & ~n3500;
  assign n3502 = n3501 ^ n3362;
  assign n3542 = n3541 ^ n3502;
  assign n3492 = n575 & n2527;
  assign n3493 = x70 & n2690;
  assign n3494 = x72 & n2693;
  assign n3495 = ~n3493 & ~n3494;
  assign n3496 = x71 & n2530;
  assign n3497 = n3495 & ~n3496;
  assign n3498 = ~n3492 & n3497;
  assign n3499 = n3498 ^ x29;
  assign n3543 = n3542 ^ n3499;
  assign n3489 = n3363 ^ n3335;
  assign n3490 = ~n3364 & ~n3489;
  assign n3491 = n3490 ^ n3335;
  assign n3544 = n3543 ^ n3491;
  assign n3481 = n789 & n2102;
  assign n3482 = x73 & n2112;
  assign n3483 = x74 & n2105;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = x75 & n2381;
  assign n3486 = n3484 & ~n3485;
  assign n3487 = ~n3481 & n3486;
  assign n3488 = n3487 ^ x26;
  assign n3545 = n3544 ^ n3488;
  assign n3478 = n3365 ^ n3324;
  assign n3479 = n3366 & n3478;
  assign n3480 = n3479 ^ n3324;
  assign n3546 = n3545 ^ n3480;
  assign n3470 = n1041 & n1746;
  assign n3471 = x76 & n1871;
  assign n3472 = x78 & n1873;
  assign n3473 = ~n3471 & ~n3472;
  assign n3474 = x77 & n1750;
  assign n3475 = n3473 & ~n3474;
  assign n3476 = ~n3470 & n3475;
  assign n3477 = n3476 ^ x23;
  assign n3547 = n3546 ^ n3477;
  assign n3467 = n3367 ^ n3313;
  assign n3468 = ~n3368 & ~n3467;
  assign n3469 = n3468 ^ n3313;
  assign n3548 = n3547 ^ n3469;
  assign n3459 = n1340 & n1404;
  assign n3460 = x79 & n1514;
  assign n3461 = x81 & n1517;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = x80 & n1408;
  assign n3464 = n3462 & ~n3463;
  assign n3465 = ~n3459 & n3464;
  assign n3466 = n3465 ^ x20;
  assign n3549 = n3548 ^ n3466;
  assign n3456 = n3369 ^ n3302;
  assign n3457 = n3370 & n3456;
  assign n3458 = n3457 ^ n3302;
  assign n3550 = n3549 ^ n3458;
  assign n3448 = n1098 & n1667;
  assign n3449 = x83 & n1102;
  assign n3450 = x82 & n1198;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = x84 & n1201;
  assign n3453 = n3451 & ~n3452;
  assign n3454 = ~n3448 & n3453;
  assign n3455 = n3454 ^ x17;
  assign n3551 = n3550 ^ n3455;
  assign n3445 = n3371 ^ n3291;
  assign n3446 = ~n3372 & ~n3445;
  assign n3447 = n3446 ^ n3291;
  assign n3552 = n3551 ^ n3447;
  assign n3437 = n821 & n2039;
  assign n3438 = x85 & n898;
  assign n3439 = x86 & n824;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = x87 & n901;
  assign n3442 = n3440 & ~n3441;
  assign n3443 = ~n3437 & n3442;
  assign n3444 = n3443 ^ x14;
  assign n3553 = n3552 ^ n3444;
  assign n3434 = n3373 ^ n3280;
  assign n3435 = n3374 & n3434;
  assign n3436 = n3435 ^ n3280;
  assign n3554 = n3553 ^ n3436;
  assign n3426 = n596 & n2448;
  assign n3427 = x88 & n673;
  assign n3428 = x90 & n676;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = x89 & n601;
  assign n3431 = n3429 & ~n3430;
  assign n3432 = ~n3426 & n3431;
  assign n3433 = n3432 ^ x11;
  assign n3555 = n3554 ^ n3433;
  assign n3423 = n3375 ^ n3269;
  assign n3424 = ~n3376 & ~n3423;
  assign n3425 = n3424 ^ n3269;
  assign n3556 = n3555 ^ n3425;
  assign n3415 = n399 & n2901;
  assign n3416 = x91 & n478;
  assign n3417 = x93 & n470;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = x92 & n402;
  assign n3420 = n3418 & ~n3419;
  assign n3421 = ~n3415 & n3420;
  assign n3422 = n3421 ^ x8;
  assign n3557 = n3556 ^ n3422;
  assign n3412 = n3377 ^ n3258;
  assign n3413 = n3378 & n3412;
  assign n3414 = n3413 ^ n3258;
  assign n3558 = n3557 ^ n3414;
  assign n3403 = n2891 ^ x96;
  assign n3404 = n239 & n3403;
  assign n3405 = x94 & n249;
  assign n3406 = x95 & n242;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = x96 & n280;
  assign n3409 = n3407 & ~n3408;
  assign n3410 = ~n3404 & n3409;
  assign n3411 = n3410 ^ x5;
  assign n3559 = n3558 ^ n3411;
  assign n3400 = n3379 ^ n3246;
  assign n3401 = ~n3380 & n3400;
  assign n3402 = n3401 ^ n3246;
  assign n3560 = n3559 ^ n3402;
  assign n3392 = x98 ^ x97;
  assign n3393 = ~n3230 & n3392;
  assign n3394 = n169 & ~n3393;
  assign n3395 = n3394 ^ x1;
  assign n3396 = n3395 ^ x99;
  assign n3388 = x2 & ~x97;
  assign n3387 = x98 ^ x2;
  assign n3389 = n3388 ^ n3387;
  assign n3390 = x1 & n3389;
  assign n3391 = n3390 ^ n3388;
  assign n3397 = n3396 ^ n3391;
  assign n3398 = ~x0 & n3397;
  assign n3399 = n3398 ^ n3396;
  assign n3561 = n3560 ^ n3399;
  assign n3384 = n3381 ^ n3216;
  assign n3385 = n3382 & ~n3384;
  assign n3386 = n3385 ^ n3216;
  assign n3562 = n3561 ^ n3386;
  assign n3710 = n3516 & n3539;
  assign n3695 = n3356 ^ x35;
  assign n3696 = n3695 ^ n3356;
  assign n3697 = n3524 & n3696;
  assign n3698 = n3697 ^ n3356;
  assign n3699 = n3521 & n3698;
  assign n3700 = x65 & n3699;
  assign n3701 = n3175 & ~n3521;
  assign n3702 = x67 & n3701;
  assign n3703 = ~n3700 & ~n3702;
  assign n3704 = x66 & n3526;
  assign n3705 = n3703 & ~n3704;
  assign n3706 = n285 & n3522;
  assign n3707 = n3705 & ~n3706;
  assign n3708 = n3707 ^ x35;
  assign n3693 = x36 ^ x35;
  assign n3694 = x64 & n3693;
  assign n3709 = n3708 ^ n3694;
  assign n3711 = n3710 ^ n3709;
  assign n3685 = n458 & n3009;
  assign n3686 = x68 & n3181;
  assign n3687 = x70 & n3183;
  assign n3688 = ~n3686 & ~n3687;
  assign n3689 = x69 & n3013;
  assign n3690 = n3688 & ~n3689;
  assign n3691 = ~n3685 & n3690;
  assign n3692 = n3691 ^ x32;
  assign n3712 = n3711 ^ n3692;
  assign n3682 = n3540 ^ n3502;
  assign n3683 = n3541 & n3682;
  assign n3684 = n3683 ^ n3502;
  assign n3713 = n3712 ^ n3684;
  assign n3674 = ~n653 & n2527;
  assign n3675 = x71 & n2690;
  assign n3676 = x73 & n2693;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = x72 & n2530;
  assign n3679 = n3677 & ~n3678;
  assign n3680 = ~n3674 & n3679;
  assign n3681 = n3680 ^ x29;
  assign n3714 = n3713 ^ n3681;
  assign n3671 = n3542 ^ n3491;
  assign n3672 = ~n3543 & ~n3671;
  assign n3673 = n3672 ^ n3491;
  assign n3715 = n3714 ^ n3673;
  assign n3663 = n870 & n2102;
  assign n3664 = x74 & n2112;
  assign n3665 = x76 & n2381;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = x75 & n2105;
  assign n3668 = n3666 & ~n3667;
  assign n3669 = ~n3663 & n3668;
  assign n3670 = n3669 ^ x26;
  assign n3716 = n3715 ^ n3670;
  assign n3660 = n3544 ^ n3480;
  assign n3661 = n3545 & n3660;
  assign n3662 = n3661 ^ n3480;
  assign n3717 = n3716 ^ n3662;
  assign n3652 = n1149 & n1746;
  assign n3653 = x77 & n1871;
  assign n3654 = x78 & n1750;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = x79 & n1873;
  assign n3657 = n3655 & ~n3656;
  assign n3658 = ~n3652 & n3657;
  assign n3659 = n3658 ^ x23;
  assign n3718 = n3717 ^ n3659;
  assign n3649 = n3546 ^ n3469;
  assign n3650 = ~n3547 & ~n3649;
  assign n3651 = n3650 ^ n3469;
  assign n3719 = n3718 ^ n3651;
  assign n3641 = n1404 & n1454;
  assign n3642 = x80 & n1514;
  assign n3643 = x81 & n1408;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = x82 & n1517;
  assign n3646 = n3644 & ~n3645;
  assign n3647 = ~n3641 & n3646;
  assign n3648 = n3647 ^ x20;
  assign n3720 = n3719 ^ n3648;
  assign n3638 = n3548 ^ n3458;
  assign n3639 = n3549 & n3638;
  assign n3640 = n3639 ^ n3458;
  assign n3721 = n3720 ^ n3640;
  assign n3630 = n1098 & n1801;
  assign n3631 = x84 & n1102;
  assign n3632 = x83 & n1198;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = x85 & n1201;
  assign n3635 = n3633 & ~n3634;
  assign n3636 = ~n3630 & n3635;
  assign n3637 = n3636 ^ x17;
  assign n3722 = n3721 ^ n3637;
  assign n3627 = n3550 ^ n3447;
  assign n3628 = ~n3551 & ~n3627;
  assign n3629 = n3628 ^ n3447;
  assign n3723 = n3722 ^ n3629;
  assign n3619 = n821 & n2176;
  assign n3620 = x86 & n898;
  assign n3621 = x87 & n824;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = x88 & n901;
  assign n3624 = n3622 & ~n3623;
  assign n3625 = ~n3619 & n3624;
  assign n3626 = n3625 ^ x14;
  assign n3724 = n3723 ^ n3626;
  assign n3616 = n3552 ^ n3436;
  assign n3617 = n3553 & n3616;
  assign n3618 = n3617 ^ n3436;
  assign n3725 = n3724 ^ n3618;
  assign n3608 = n596 & n2607;
  assign n3609 = x89 & n673;
  assign n3610 = x90 & n601;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = x91 & n676;
  assign n3613 = n3611 & ~n3612;
  assign n3614 = ~n3608 & n3613;
  assign n3615 = n3614 ^ x11;
  assign n3726 = n3725 ^ n3615;
  assign n3605 = n3554 ^ n3425;
  assign n3606 = ~n3555 & ~n3605;
  assign n3607 = n3606 ^ n3425;
  assign n3727 = n3726 ^ n3607;
  assign n3597 = n399 & n3078;
  assign n3598 = x92 & n478;
  assign n3599 = x93 & n402;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = x94 & n470;
  assign n3602 = n3600 & ~n3601;
  assign n3603 = ~n3597 & n3602;
  assign n3604 = n3603 ^ x8;
  assign n3728 = n3727 ^ n3604;
  assign n3594 = n3556 ^ n3414;
  assign n3595 = n3557 & n3594;
  assign n3596 = n3595 ^ n3414;
  assign n3729 = n3728 ^ n3596;
  assign n3585 = n3068 ^ x97;
  assign n3586 = n239 & n3585;
  assign n3587 = x95 & n249;
  assign n3588 = x97 & n280;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = x96 & n242;
  assign n3591 = n3589 & ~n3590;
  assign n3592 = ~n3586 & n3591;
  assign n3593 = n3592 ^ x5;
  assign n3730 = n3729 ^ n3593;
  assign n3582 = n3558 ^ n3402;
  assign n3583 = ~n3559 & n3582;
  assign n3584 = n3583 ^ n3402;
  assign n3731 = n3730 ^ n3584;
  assign n3568 = x99 ^ x98;
  assign n3569 = ~n3393 & n3568;
  assign n3570 = n169 & ~n3569;
  assign n3571 = n3570 ^ x1;
  assign n3572 = n3571 ^ x100;
  assign n3566 = x99 ^ x2;
  assign n3567 = x1 & n3566;
  assign n3573 = n3572 ^ n3567;
  assign n3574 = n3573 ^ n3572;
  assign n3575 = ~x98 & n197;
  assign n3576 = n3575 ^ n3572;
  assign n3577 = n3576 ^ n3572;
  assign n3578 = ~n3574 & ~n3577;
  assign n3579 = n3578 ^ n3572;
  assign n3580 = ~x0 & ~n3579;
  assign n3581 = n3580 ^ n3572;
  assign n3732 = n3731 ^ n3581;
  assign n3563 = n3560 ^ n3386;
  assign n3564 = n3561 & ~n3563;
  assign n3565 = n3564 ^ n3386;
  assign n3733 = n3732 ^ n3565;
  assign n3887 = ~n3694 & ~n3710;
  assign n3888 = ~n3708 & ~n3887;
  assign n3882 = x65 ^ x36;
  assign n3883 = n3693 & ~n3882;
  assign n3884 = n3883 ^ x35;
  assign n3885 = n3884 ^ x37;
  assign n3879 = x35 & x36;
  assign n3880 = n3879 ^ x37;
  assign n3881 = ~x64 & n3880;
  assign n3886 = n3885 ^ n3881;
  assign n3889 = n3888 ^ n3886;
  assign n3871 = n321 & n3522;
  assign n3872 = x66 & n3699;
  assign n3873 = x68 & n3701;
  assign n3874 = ~n3872 & ~n3873;
  assign n3875 = x67 & n3526;
  assign n3876 = n3874 & ~n3875;
  assign n3877 = ~n3871 & n3876;
  assign n3878 = n3877 ^ x35;
  assign n3890 = n3889 ^ n3878;
  assign n3863 = n517 & n3009;
  assign n3864 = x70 & n3013;
  assign n3865 = x69 & n3181;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = x71 & n3183;
  assign n3868 = n3866 & ~n3867;
  assign n3869 = ~n3863 & n3868;
  assign n3870 = n3869 ^ x32;
  assign n3891 = n3890 ^ n3870;
  assign n3860 = n3711 ^ n3684;
  assign n3861 = ~n3712 & ~n3860;
  assign n3862 = n3861 ^ n3684;
  assign n3892 = n3891 ^ n3862;
  assign n3852 = ~n721 & n2527;
  assign n3853 = x72 & n2690;
  assign n3854 = x74 & n2693;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = x73 & n2530;
  assign n3857 = n3855 & ~n3856;
  assign n3858 = ~n3852 & n3857;
  assign n3859 = n3858 ^ x29;
  assign n3893 = n3892 ^ n3859;
  assign n3849 = n3681 ^ n3673;
  assign n3850 = ~n3714 & n3849;
  assign n3851 = n3850 ^ n3713;
  assign n3894 = n3893 ^ n3851;
  assign n3841 = n956 & n2102;
  assign n3842 = x75 & n2112;
  assign n3843 = x77 & n2381;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = x76 & n2105;
  assign n3846 = n3844 & ~n3845;
  assign n3847 = ~n3841 & n3846;
  assign n3848 = n3847 ^ x26;
  assign n3895 = n3894 ^ n3848;
  assign n3838 = n3715 ^ n3662;
  assign n3839 = ~n3716 & ~n3838;
  assign n3840 = n3839 ^ n3662;
  assign n3896 = n3895 ^ n3840;
  assign n3830 = n1242 & n1746;
  assign n3831 = x78 & n1871;
  assign n3832 = x79 & n1750;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = x80 & n1873;
  assign n3835 = n3833 & ~n3834;
  assign n3836 = ~n3830 & n3835;
  assign n3837 = n3836 ^ x23;
  assign n3897 = n3896 ^ n3837;
  assign n3827 = n3717 ^ n3651;
  assign n3828 = n3718 & n3827;
  assign n3829 = n3828 ^ n3651;
  assign n3898 = n3897 ^ n3829;
  assign n3819 = n1404 & n1560;
  assign n3820 = x81 & n1514;
  assign n3821 = x82 & n1408;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = x83 & n1517;
  assign n3824 = n3822 & ~n3823;
  assign n3825 = ~n3819 & n3824;
  assign n3826 = n3825 ^ x20;
  assign n3899 = n3898 ^ n3826;
  assign n3816 = n3719 ^ n3640;
  assign n3817 = ~n3720 & ~n3816;
  assign n3818 = n3817 ^ n3640;
  assign n3900 = n3899 ^ n3818;
  assign n3808 = n1098 & n1920;
  assign n3809 = x85 & n1102;
  assign n3810 = x84 & n1198;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = x86 & n1201;
  assign n3813 = n3811 & ~n3812;
  assign n3814 = ~n3808 & n3813;
  assign n3815 = n3814 ^ x17;
  assign n3901 = n3900 ^ n3815;
  assign n3805 = n3721 ^ n3629;
  assign n3806 = n3722 & n3805;
  assign n3807 = n3806 ^ n3629;
  assign n3902 = n3901 ^ n3807;
  assign n3797 = n821 & n2310;
  assign n3798 = x87 & n898;
  assign n3799 = x89 & n901;
  assign n3800 = ~n3798 & ~n3799;
  assign n3801 = x88 & n824;
  assign n3802 = n3800 & ~n3801;
  assign n3803 = ~n3797 & n3802;
  assign n3804 = n3803 ^ x14;
  assign n3903 = n3902 ^ n3804;
  assign n3794 = n3723 ^ n3618;
  assign n3795 = ~n3724 & ~n3794;
  assign n3796 = n3795 ^ n3618;
  assign n3904 = n3903 ^ n3796;
  assign n3786 = n596 & n2755;
  assign n3787 = x90 & n673;
  assign n3788 = x92 & n676;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = x91 & n601;
  assign n3791 = n3789 & ~n3790;
  assign n3792 = ~n3786 & n3791;
  assign n3793 = n3792 ^ x11;
  assign n3905 = n3904 ^ n3793;
  assign n3783 = n3725 ^ n3607;
  assign n3784 = n3726 & n3783;
  assign n3785 = n3784 ^ n3607;
  assign n3906 = n3905 ^ n3785;
  assign n3775 = n399 & n3247;
  assign n3776 = x93 & n478;
  assign n3777 = x94 & n402;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = x95 & n470;
  assign n3780 = n3778 & ~n3779;
  assign n3781 = ~n3775 & n3780;
  assign n3782 = n3781 ^ x8;
  assign n3907 = n3906 ^ n3782;
  assign n3772 = n3727 ^ n3596;
  assign n3773 = ~n3728 & ~n3772;
  assign n3774 = n3773 ^ n3596;
  assign n3908 = n3907 ^ n3774;
  assign n3763 = n3392 ^ n3229;
  assign n3764 = n239 & n3763;
  assign n3765 = x96 & n249;
  assign n3766 = x98 & n280;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = x97 & n242;
  assign n3769 = n3767 & ~n3768;
  assign n3770 = ~n3764 & n3769;
  assign n3771 = n3770 ^ x5;
  assign n3909 = n3908 ^ n3771;
  assign n3760 = n3729 ^ n3584;
  assign n3761 = n3730 & ~n3760;
  assign n3762 = n3761 ^ n3584;
  assign n3910 = n3909 ^ n3762;
  assign n3749 = x100 ^ x99;
  assign n3750 = x100 ^ x98;
  assign n3751 = ~n3393 & ~n3750;
  assign n3752 = n3749 & n3751;
  assign n3753 = n3752 ^ n3749;
  assign n3754 = n169 & ~n3753;
  assign n3755 = n3754 ^ x1;
  assign n3756 = n3755 ^ x101;
  assign n3737 = x100 ^ x2;
  assign n3738 = n3737 ^ x1;
  assign n3739 = n3738 ^ n3737;
  assign n3740 = n3739 ^ x0;
  assign n3741 = n3737 ^ x100;
  assign n3742 = n3741 ^ x99;
  assign n3743 = ~x99 & ~n3742;
  assign n3744 = n3743 ^ n3737;
  assign n3745 = n3744 ^ x99;
  assign n3746 = n3740 & ~n3745;
  assign n3747 = n3746 ^ n3743;
  assign n3748 = n3747 ^ x99;
  assign n3757 = n3756 ^ n3748;
  assign n3758 = ~x0 & ~n3757;
  assign n3759 = n3758 ^ n3756;
  assign n3911 = n3910 ^ n3759;
  assign n3734 = n3731 ^ n3565;
  assign n3735 = ~n3732 & n3734;
  assign n3736 = n3735 ^ n3565;
  assign n3912 = n3911 ^ n3736;
  assign n4092 = n1340 & n1746;
  assign n4093 = x80 & n1750;
  assign n4094 = x79 & n1871;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = x81 & n1873;
  assign n4097 = n4095 & ~n4096;
  assign n4098 = ~n4092 & n4097;
  assign n4099 = n4098 ^ x23;
  assign n4089 = n3896 ^ n3829;
  assign n4090 = n3897 & n4089;
  assign n4091 = n4090 ^ n3829;
  assign n4100 = n4099 ^ n4091;
  assign n4079 = n1041 & n2102;
  assign n4080 = x76 & n2112;
  assign n4081 = x77 & n2105;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = x78 & n2381;
  assign n4084 = n4082 & ~n4083;
  assign n4085 = ~n4079 & n4084;
  assign n4086 = n4085 ^ x26;
  assign n4076 = n3894 ^ n3840;
  assign n4077 = ~n3895 & ~n4076;
  assign n4078 = n4077 ^ n3840;
  assign n4087 = n4086 ^ n4078;
  assign n4066 = n789 & n2527;
  assign n4067 = x74 & n2530;
  assign n4068 = x73 & n2690;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = x75 & n2693;
  assign n4071 = n4069 & ~n4070;
  assign n4072 = ~n4066 & n4071;
  assign n4073 = n4072 ^ x29;
  assign n4063 = n3892 ^ n3851;
  assign n4064 = n3893 & n4063;
  assign n4065 = n4064 ^ n3851;
  assign n4074 = n4073 ^ n4065;
  assign n4035 = ~x35 & ~x36;
  assign n4036 = ~x37 & x38;
  assign n4037 = n4035 & n4036;
  assign n4038 = x64 & n4037;
  assign n4039 = x38 ^ x37;
  assign n4040 = n3693 & n4039;
  assign n4041 = n142 & n4040;
  assign n4042 = n4035 ^ n3879;
  assign n4043 = x37 & n4042;
  assign n4044 = n4043 ^ n3879;
  assign n4045 = ~n4041 & ~n4044;
  assign n4046 = x65 & ~n4045;
  assign n4047 = n152 & n4039;
  assign n4048 = x66 & n3693;
  assign n4049 = ~n4047 & n4048;
  assign n4050 = ~n4046 & ~n4049;
  assign n4051 = n4050 ^ x38;
  assign n4052 = x37 & x64;
  assign n4053 = n3879 & n4052;
  assign n4054 = n4050 & n4053;
  assign n4055 = n4051 & n4054;
  assign n4056 = n4055 ^ n4051;
  assign n4057 = ~n4038 & ~n4056;
  assign n4029 = x37 ^ x35;
  assign n4030 = x64 & n4029;
  assign n4031 = n4030 ^ n233;
  assign n4032 = ~n3693 & ~n4031;
  assign n4033 = n4032 ^ n233;
  assign n4034 = x38 & n4033;
  assign n4058 = n4057 ^ n4034;
  assign n4021 = n420 & n3522;
  assign n4022 = x68 & n3526;
  assign n4023 = x67 & n3699;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = x69 & n3701;
  assign n4026 = n4024 & ~n4025;
  assign n4027 = ~n4021 & n4026;
  assign n4028 = n4027 ^ x35;
  assign n4059 = n4058 ^ n4028;
  assign n4018 = n3886 ^ n3878;
  assign n4019 = n3889 & n4018;
  assign n4020 = n4019 ^ n3888;
  assign n4060 = n4059 ^ n4020;
  assign n4010 = n575 & n3009;
  assign n4011 = x70 & n3181;
  assign n4012 = x72 & n3183;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = x71 & n3013;
  assign n4015 = n4013 & ~n4014;
  assign n4016 = ~n4010 & n4015;
  assign n4017 = n4016 ^ x32;
  assign n4061 = n4060 ^ n4017;
  assign n4007 = n3890 ^ n3862;
  assign n4008 = ~n3891 & ~n4007;
  assign n4009 = n4008 ^ n3862;
  assign n4062 = n4061 ^ n4009;
  assign n4075 = n4074 ^ n4062;
  assign n4088 = n4087 ^ n4075;
  assign n4101 = n4100 ^ n4088;
  assign n3999 = n1404 & n1667;
  assign n4000 = x82 & n1514;
  assign n4001 = x83 & n1408;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = x84 & n1517;
  assign n4004 = n4002 & ~n4003;
  assign n4005 = ~n3999 & n4004;
  assign n4006 = n4005 ^ x20;
  assign n4102 = n4101 ^ n4006;
  assign n3996 = n3898 ^ n3818;
  assign n3997 = ~n3899 & ~n3996;
  assign n3998 = n3997 ^ n3818;
  assign n4103 = n4102 ^ n3998;
  assign n3988 = n1098 & n2039;
  assign n3989 = x86 & n1102;
  assign n3990 = x85 & n1198;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = x87 & n1201;
  assign n3993 = n3991 & ~n3992;
  assign n3994 = ~n3988 & n3993;
  assign n3995 = n3994 ^ x17;
  assign n4104 = n4103 ^ n3995;
  assign n3985 = n3900 ^ n3807;
  assign n3986 = n3901 & n3985;
  assign n3987 = n3986 ^ n3807;
  assign n4105 = n4104 ^ n3987;
  assign n3977 = n821 & n2448;
  assign n3978 = x88 & n898;
  assign n3979 = x90 & n901;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = x89 & n824;
  assign n3982 = n3980 & ~n3981;
  assign n3983 = ~n3977 & n3982;
  assign n3984 = n3983 ^ x14;
  assign n4106 = n4105 ^ n3984;
  assign n3974 = n3902 ^ n3796;
  assign n3975 = ~n3903 & ~n3974;
  assign n3976 = n3975 ^ n3796;
  assign n4107 = n4106 ^ n3976;
  assign n3966 = n596 & n2901;
  assign n3967 = x91 & n673;
  assign n3968 = x92 & n601;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = x93 & n676;
  assign n3971 = n3969 & ~n3970;
  assign n3972 = ~n3966 & n3971;
  assign n3973 = n3972 ^ x11;
  assign n4108 = n4107 ^ n3973;
  assign n3963 = n3904 ^ n3785;
  assign n3964 = n3905 & n3963;
  assign n3965 = n3964 ^ n3785;
  assign n4109 = n4108 ^ n3965;
  assign n3955 = n399 & n3403;
  assign n3956 = x94 & n478;
  assign n3957 = x95 & n402;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = x96 & n470;
  assign n3960 = n3958 & ~n3959;
  assign n3961 = ~n3955 & n3960;
  assign n3962 = n3961 ^ x8;
  assign n4110 = n4109 ^ n3962;
  assign n3952 = n3906 ^ n3774;
  assign n3953 = ~n3907 & ~n3952;
  assign n3954 = n3953 ^ n3774;
  assign n4111 = n4110 ^ n3954;
  assign n3943 = n3393 ^ x99;
  assign n3944 = n239 & n3943;
  assign n3945 = x98 & n242;
  assign n3946 = x97 & n249;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = x99 & n280;
  assign n3949 = n3947 & ~n3948;
  assign n3950 = ~n3944 & n3949;
  assign n3951 = n3950 ^ x5;
  assign n4112 = n4111 ^ n3951;
  assign n3940 = n3908 ^ n3762;
  assign n3941 = n3909 & ~n3940;
  assign n3942 = n3941 ^ n3762;
  assign n4113 = n4112 ^ n3942;
  assign n3925 = ~x98 & ~n3393;
  assign n3926 = x99 & x101;
  assign n3927 = ~n3925 & n3926;
  assign n3928 = ~x100 & ~n3927;
  assign n3929 = x98 & ~n3393;
  assign n3930 = ~x99 & ~x101;
  assign n3931 = ~n3929 & n3930;
  assign n3932 = ~n3928 & ~n3931;
  assign n3933 = n3932 ^ x101;
  assign n3934 = n169 & ~n3933;
  assign n3935 = n3934 ^ x1;
  assign n3936 = n3935 ^ x102;
  assign n3916 = x101 ^ x2;
  assign n3917 = n3916 ^ x101;
  assign n3918 = x101 ^ x100;
  assign n3919 = n3918 ^ x101;
  assign n3920 = n3917 & n3919;
  assign n3921 = n3920 ^ x101;
  assign n3922 = ~x1 & n3921;
  assign n3923 = n3922 ^ x101;
  assign n3924 = n3923 ^ x2;
  assign n3937 = n3936 ^ n3924;
  assign n3938 = ~x0 & n3937;
  assign n3939 = n3938 ^ n3936;
  assign n4114 = n4113 ^ n3939;
  assign n3913 = n3910 ^ n3736;
  assign n3914 = ~n3911 & n3913;
  assign n3915 = n3914 ^ n3736;
  assign n4115 = n4114 ^ n3915;
  assign n4277 = n4034 & n4057;
  assign n4262 = x66 & n4044;
  assign n4263 = n3879 ^ x38;
  assign n4264 = n4263 ^ n3879;
  assign n4265 = n4042 & n4264;
  assign n4266 = n4265 ^ n3879;
  assign n4267 = n4039 & n4266;
  assign n4268 = x65 & n4267;
  assign n4269 = ~n4262 & ~n4268;
  assign n4270 = n3693 & ~n4039;
  assign n4271 = x67 & n4270;
  assign n4272 = n4269 & ~n4271;
  assign n4273 = n285 & n4040;
  assign n4274 = n4272 & ~n4273;
  assign n4275 = n4274 ^ x38;
  assign n4260 = x39 ^ x38;
  assign n4261 = x64 & n4260;
  assign n4276 = n4275 ^ n4261;
  assign n4278 = n4277 ^ n4276;
  assign n4252 = n458 & n3522;
  assign n4253 = x68 & n3699;
  assign n4254 = x69 & n3526;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = x70 & n3701;
  assign n4257 = n4255 & ~n4256;
  assign n4258 = ~n4252 & n4257;
  assign n4259 = n4258 ^ x35;
  assign n4279 = n4278 ^ n4259;
  assign n4249 = n4058 ^ n4020;
  assign n4250 = n4059 & n4249;
  assign n4251 = n4250 ^ n4020;
  assign n4280 = n4279 ^ n4251;
  assign n4241 = ~n653 & n3009;
  assign n4242 = x72 & n3013;
  assign n4243 = x73 & n3183;
  assign n4244 = ~n4242 & ~n4243;
  assign n4245 = x71 & n3181;
  assign n4246 = n4244 & ~n4245;
  assign n4247 = ~n4241 & n4246;
  assign n4248 = n4247 ^ x32;
  assign n4281 = n4280 ^ n4248;
  assign n4238 = n4060 ^ n4009;
  assign n4239 = ~n4061 & ~n4238;
  assign n4240 = n4239 ^ n4009;
  assign n4282 = n4281 ^ n4240;
  assign n4230 = n870 & n2527;
  assign n4231 = x74 & n2690;
  assign n4232 = x76 & n2693;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = x75 & n2530;
  assign n4235 = n4233 & ~n4234;
  assign n4236 = ~n4230 & n4235;
  assign n4237 = n4236 ^ x29;
  assign n4283 = n4282 ^ n4237;
  assign n4227 = n4073 ^ n4062;
  assign n4228 = ~n4074 & n4227;
  assign n4229 = n4228 ^ n4065;
  assign n4284 = n4283 ^ n4229;
  assign n4219 = n1149 & n2102;
  assign n4220 = x77 & n2112;
  assign n4221 = x79 & n2381;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = x78 & n2105;
  assign n4224 = n4222 & ~n4223;
  assign n4225 = ~n4219 & n4224;
  assign n4226 = n4225 ^ x26;
  assign n4285 = n4284 ^ n4226;
  assign n4216 = n4086 ^ n4075;
  assign n4217 = ~n4087 & ~n4216;
  assign n4218 = n4217 ^ n4078;
  assign n4286 = n4285 ^ n4218;
  assign n4208 = n1454 & n1746;
  assign n4209 = x80 & n1871;
  assign n4210 = x81 & n1750;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = x82 & n1873;
  assign n4213 = n4211 & ~n4212;
  assign n4214 = ~n4208 & n4213;
  assign n4215 = n4214 ^ x23;
  assign n4287 = n4286 ^ n4215;
  assign n4205 = n4099 ^ n4088;
  assign n4206 = ~n4100 & n4205;
  assign n4207 = n4206 ^ n4091;
  assign n4288 = n4287 ^ n4207;
  assign n4197 = n1404 & n1801;
  assign n4198 = x83 & n1514;
  assign n4199 = x84 & n1408;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = x85 & n1517;
  assign n4202 = n4200 & ~n4201;
  assign n4203 = ~n4197 & n4202;
  assign n4204 = n4203 ^ x20;
  assign n4289 = n4288 ^ n4204;
  assign n4194 = n4101 ^ n3998;
  assign n4195 = ~n4102 & ~n4194;
  assign n4196 = n4195 ^ n3998;
  assign n4290 = n4289 ^ n4196;
  assign n4186 = n1098 & n2176;
  assign n4187 = x87 & n1102;
  assign n4188 = x86 & n1198;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = x88 & n1201;
  assign n4191 = n4189 & ~n4190;
  assign n4192 = ~n4186 & n4191;
  assign n4193 = n4192 ^ x17;
  assign n4291 = n4290 ^ n4193;
  assign n4183 = n4103 ^ n3987;
  assign n4184 = n4104 & n4183;
  assign n4185 = n4184 ^ n3987;
  assign n4292 = n4291 ^ n4185;
  assign n4175 = n821 & n2607;
  assign n4176 = x89 & n898;
  assign n4177 = x91 & n901;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = x90 & n824;
  assign n4180 = n4178 & ~n4179;
  assign n4181 = ~n4175 & n4180;
  assign n4182 = n4181 ^ x14;
  assign n4293 = n4292 ^ n4182;
  assign n4172 = n4105 ^ n3976;
  assign n4173 = ~n4106 & ~n4172;
  assign n4174 = n4173 ^ n3976;
  assign n4294 = n4293 ^ n4174;
  assign n4164 = n596 & n3078;
  assign n4165 = x92 & n673;
  assign n4166 = x94 & n676;
  assign n4167 = ~n4165 & ~n4166;
  assign n4168 = x93 & n601;
  assign n4169 = n4167 & ~n4168;
  assign n4170 = ~n4164 & n4169;
  assign n4171 = n4170 ^ x11;
  assign n4295 = n4294 ^ n4171;
  assign n4161 = n4107 ^ n3965;
  assign n4162 = n4108 & n4161;
  assign n4163 = n4162 ^ n3965;
  assign n4296 = n4295 ^ n4163;
  assign n4153 = n399 & n3585;
  assign n4154 = x95 & n478;
  assign n4155 = x97 & n470;
  assign n4156 = ~n4154 & ~n4155;
  assign n4157 = x96 & n402;
  assign n4158 = n4156 & ~n4157;
  assign n4159 = ~n4153 & n4158;
  assign n4160 = n4159 ^ x8;
  assign n4297 = n4296 ^ n4160;
  assign n4150 = n4109 ^ n3954;
  assign n4151 = ~n4110 & ~n4150;
  assign n4152 = n4151 ^ n3954;
  assign n4298 = n4297 ^ n4152;
  assign n4141 = n3569 ^ x100;
  assign n4142 = n239 & n4141;
  assign n4143 = x98 & n249;
  assign n4144 = x99 & n242;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = x100 & n280;
  assign n4147 = n4145 & ~n4146;
  assign n4148 = ~n4142 & n4147;
  assign n4149 = n4148 ^ x5;
  assign n4299 = n4298 ^ n4149;
  assign n4138 = n4111 ^ n3942;
  assign n4139 = n4112 & ~n4138;
  assign n4140 = n4139 ^ n3942;
  assign n4300 = n4299 ^ n4140;
  assign n4127 = x101 & n3932;
  assign n4128 = ~x102 & ~n4127;
  assign n4129 = ~x101 & ~n3932;
  assign n4130 = x102 & ~n4129;
  assign n4131 = ~n4128 & ~n4130;
  assign n4132 = n169 & ~n4131;
  assign n4133 = n4132 ^ x1;
  assign n4134 = n4133 ^ x103;
  assign n4119 = x102 ^ x2;
  assign n4120 = n4119 ^ x101;
  assign n4121 = n4120 ^ n4119;
  assign n4122 = n4119 ^ x102;
  assign n4123 = ~n4121 & n4122;
  assign n4124 = n4123 ^ n4119;
  assign n4125 = ~x1 & n4124;
  assign n4126 = n4125 ^ n4119;
  assign n4135 = n4134 ^ n4126;
  assign n4136 = ~x0 & n4135;
  assign n4137 = n4136 ^ n4134;
  assign n4301 = n4300 ^ n4137;
  assign n4116 = n4113 ^ n3915;
  assign n4117 = ~n4114 & n4116;
  assign n4118 = n4117 ^ n3915;
  assign n4302 = n4301 ^ n4118;
  assign n4454 = n517 & n3522;
  assign n4455 = x70 & n3526;
  assign n4456 = x69 & n3699;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = x71 & n3701;
  assign n4459 = n4457 & ~n4458;
  assign n4460 = ~n4454 & n4459;
  assign n4461 = n4460 ^ x35;
  assign n4451 = n4278 ^ n4251;
  assign n4452 = ~n4279 & ~n4451;
  assign n4453 = n4452 ^ n4251;
  assign n4462 = n4461 ^ n4453;
  assign n4445 = x38 & x39;
  assign n4446 = n4445 ^ x40;
  assign n4447 = ~x64 & n4446;
  assign n4441 = x65 ^ x39;
  assign n4442 = n4260 & ~n4441;
  assign n4443 = n4442 ^ x38;
  assign n4444 = n4443 ^ x40;
  assign n4448 = n4447 ^ n4444;
  assign n4439 = ~n4261 & ~n4277;
  assign n4440 = ~n4275 & ~n4439;
  assign n4449 = n4448 ^ n4440;
  assign n4431 = n321 & n4040;
  assign n4432 = x67 & n4044;
  assign n4433 = x66 & n4267;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = x68 & n4270;
  assign n4436 = n4434 & ~n4435;
  assign n4437 = ~n4431 & n4436;
  assign n4438 = n4437 ^ x38;
  assign n4450 = n4449 ^ n4438;
  assign n4463 = n4462 ^ n4450;
  assign n4423 = ~n721 & n3009;
  assign n4424 = x72 & n3181;
  assign n4425 = x74 & n3183;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = x73 & n3013;
  assign n4428 = n4426 & ~n4427;
  assign n4429 = ~n4423 & n4428;
  assign n4430 = n4429 ^ x32;
  assign n4464 = n4463 ^ n4430;
  assign n4420 = n4280 ^ n4240;
  assign n4421 = n4281 & n4420;
  assign n4422 = n4421 ^ n4240;
  assign n4465 = n4464 ^ n4422;
  assign n4412 = n956 & n2527;
  assign n4413 = x76 & n2530;
  assign n4414 = x75 & n2690;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = x77 & n2693;
  assign n4417 = n4415 & ~n4416;
  assign n4418 = ~n4412 & n4417;
  assign n4419 = n4418 ^ x29;
  assign n4466 = n4465 ^ n4419;
  assign n4409 = n4282 ^ n4229;
  assign n4410 = ~n4283 & ~n4409;
  assign n4411 = n4410 ^ n4229;
  assign n4467 = n4466 ^ n4411;
  assign n4401 = n1242 & n2102;
  assign n4402 = x79 & n2105;
  assign n4403 = x80 & n2381;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = x78 & n2112;
  assign n4406 = n4404 & ~n4405;
  assign n4407 = ~n4401 & n4406;
  assign n4408 = n4407 ^ x26;
  assign n4468 = n4467 ^ n4408;
  assign n4398 = n4284 ^ n4218;
  assign n4399 = n4285 & n4398;
  assign n4400 = n4399 ^ n4218;
  assign n4469 = n4468 ^ n4400;
  assign n4390 = n1560 & n1746;
  assign n4391 = x81 & n1871;
  assign n4392 = x82 & n1750;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = x83 & n1873;
  assign n4395 = n4393 & ~n4394;
  assign n4396 = ~n4390 & n4395;
  assign n4397 = n4396 ^ x23;
  assign n4470 = n4469 ^ n4397;
  assign n4387 = n4286 ^ n4207;
  assign n4388 = ~n4287 & ~n4387;
  assign n4389 = n4388 ^ n4207;
  assign n4471 = n4470 ^ n4389;
  assign n4379 = n1404 & n1920;
  assign n4380 = x84 & n1514;
  assign n4381 = x86 & n1517;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = x85 & n1408;
  assign n4384 = n4382 & ~n4383;
  assign n4385 = ~n4379 & n4384;
  assign n4386 = n4385 ^ x20;
  assign n4472 = n4471 ^ n4386;
  assign n4376 = n4288 ^ n4196;
  assign n4377 = n4289 & n4376;
  assign n4378 = n4377 ^ n4196;
  assign n4473 = n4472 ^ n4378;
  assign n4368 = n1098 & n2310;
  assign n4369 = x88 & n1102;
  assign n4370 = x87 & n1198;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = x89 & n1201;
  assign n4373 = n4371 & ~n4372;
  assign n4374 = ~n4368 & n4373;
  assign n4375 = n4374 ^ x17;
  assign n4474 = n4473 ^ n4375;
  assign n4365 = n4290 ^ n4185;
  assign n4366 = ~n4291 & ~n4365;
  assign n4367 = n4366 ^ n4185;
  assign n4475 = n4474 ^ n4367;
  assign n4357 = n821 & n2755;
  assign n4358 = x90 & n898;
  assign n4359 = x91 & n824;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = x92 & n901;
  assign n4362 = n4360 & ~n4361;
  assign n4363 = ~n4357 & n4362;
  assign n4364 = n4363 ^ x14;
  assign n4476 = n4475 ^ n4364;
  assign n4354 = n4292 ^ n4174;
  assign n4355 = n4293 & n4354;
  assign n4356 = n4355 ^ n4174;
  assign n4477 = n4476 ^ n4356;
  assign n4346 = n596 & n3247;
  assign n4347 = x93 & n673;
  assign n4348 = x95 & n676;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = x94 & n601;
  assign n4351 = n4349 & ~n4350;
  assign n4352 = ~n4346 & n4351;
  assign n4353 = n4352 ^ x11;
  assign n4478 = n4477 ^ n4353;
  assign n4343 = n4294 ^ n4163;
  assign n4344 = ~n4295 & ~n4343;
  assign n4345 = n4344 ^ n4163;
  assign n4479 = n4478 ^ n4345;
  assign n4335 = n399 & n3763;
  assign n4336 = x96 & n478;
  assign n4337 = x98 & n470;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = x97 & n402;
  assign n4340 = n4338 & ~n4339;
  assign n4341 = ~n4335 & n4340;
  assign n4342 = n4341 ^ x8;
  assign n4480 = n4479 ^ n4342;
  assign n4332 = n4296 ^ n4152;
  assign n4333 = n4297 & n4332;
  assign n4334 = n4333 ^ n4152;
  assign n4481 = n4480 ^ n4334;
  assign n4323 = n3753 ^ x101;
  assign n4324 = n239 & n4323;
  assign n4325 = x99 & n249;
  assign n4326 = x100 & n242;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = x101 & n280;
  assign n4329 = n4327 & ~n4328;
  assign n4330 = ~n4324 & n4329;
  assign n4331 = n4330 ^ x5;
  assign n4482 = n4481 ^ n4331;
  assign n4320 = n4298 ^ n4140;
  assign n4321 = ~n4299 & n4320;
  assign n4322 = n4321 ^ n4140;
  assign n4483 = n4482 ^ n4322;
  assign n4311 = x103 & ~n4128;
  assign n4312 = ~x103 & ~n4130;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = n169 & ~n4313;
  assign n4315 = n4314 ^ x1;
  assign n4316 = n4315 ^ x104;
  assign n4307 = x103 ^ x2;
  assign n4306 = x2 & ~x102;
  assign n4308 = n4307 ^ n4306;
  assign n4309 = ~x1 & n4308;
  assign n4310 = n4309 ^ n4307;
  assign n4317 = n4316 ^ n4310;
  assign n4318 = ~x0 & n4317;
  assign n4319 = n4318 ^ n4316;
  assign n4484 = n4483 ^ n4319;
  assign n4303 = n4300 ^ n4118;
  assign n4304 = n4301 & ~n4303;
  assign n4305 = n4304 ^ n4118;
  assign n4485 = n4484 ^ n4305;
  assign n4661 = n420 & n4040;
  assign n4662 = x68 & n4044;
  assign n4663 = x67 & n4267;
  assign n4664 = ~n4662 & ~n4663;
  assign n4665 = x69 & n4270;
  assign n4666 = n4664 & ~n4665;
  assign n4667 = ~n4661 & n4666;
  assign n4668 = n4667 ^ x38;
  assign n4642 = x41 ^ x40;
  assign n4643 = n4260 & n4642;
  assign n4644 = n142 & n4643;
  assign n4632 = ~x38 & ~x39;
  assign n4633 = n4632 ^ n4445;
  assign n4645 = x40 & n4633;
  assign n4646 = n4645 ^ n4445;
  assign n4647 = ~n4644 & ~n4646;
  assign n4648 = x65 & ~n4647;
  assign n4649 = n4445 ^ x41;
  assign n4650 = n4649 ^ n4445;
  assign n4651 = n4633 & n4650;
  assign n4652 = n4651 ^ n4445;
  assign n4653 = n4642 & n4652;
  assign n4654 = x64 & n4653;
  assign n4655 = n152 & n4642;
  assign n4656 = x66 & n4260;
  assign n4657 = ~n4655 & n4656;
  assign n4658 = ~n4654 & ~n4657;
  assign n4659 = ~n4648 & n4658;
  assign n4631 = x41 & ~n233;
  assign n4634 = n4632 ^ x40;
  assign n4635 = x64 ^ x40;
  assign n4636 = n4635 ^ x40;
  assign n4637 = ~n4634 & ~n4636;
  assign n4638 = n4637 ^ x40;
  assign n4639 = n4633 & ~n4638;
  assign n4640 = n4639 ^ n4445;
  assign n4641 = n4631 & ~n4640;
  assign n4660 = n4659 ^ n4641;
  assign n4669 = n4668 ^ n4660;
  assign n4628 = n4448 ^ n4438;
  assign n4629 = n4449 & n4628;
  assign n4630 = n4629 ^ n4440;
  assign n4670 = n4669 ^ n4630;
  assign n4620 = n575 & n3522;
  assign n4621 = x71 & n3526;
  assign n4622 = x72 & n3701;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = x70 & n3699;
  assign n4625 = n4623 & ~n4624;
  assign n4626 = ~n4620 & n4625;
  assign n4627 = n4626 ^ x35;
  assign n4671 = n4670 ^ n4627;
  assign n4617 = n4461 ^ n4450;
  assign n4618 = ~n4462 & ~n4617;
  assign n4619 = n4618 ^ n4453;
  assign n4672 = n4671 ^ n4619;
  assign n4609 = n789 & n3009;
  assign n4610 = x73 & n3181;
  assign n4611 = x74 & n3013;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = x75 & n3183;
  assign n4614 = n4612 & ~n4613;
  assign n4615 = ~n4609 & n4614;
  assign n4616 = n4615 ^ x32;
  assign n4673 = n4672 ^ n4616;
  assign n4606 = n4463 ^ n4422;
  assign n4607 = n4464 & n4606;
  assign n4608 = n4607 ^ n4422;
  assign n4674 = n4673 ^ n4608;
  assign n4598 = n1041 & n2527;
  assign n4599 = x76 & n2690;
  assign n4600 = x78 & n2693;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = x77 & n2530;
  assign n4603 = n4601 & ~n4602;
  assign n4604 = ~n4598 & n4603;
  assign n4605 = n4604 ^ x29;
  assign n4675 = n4674 ^ n4605;
  assign n4595 = n4465 ^ n4411;
  assign n4596 = ~n4466 & ~n4595;
  assign n4597 = n4596 ^ n4411;
  assign n4676 = n4675 ^ n4597;
  assign n4587 = n1340 & n2102;
  assign n4588 = x79 & n2112;
  assign n4589 = x81 & n2381;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = x80 & n2105;
  assign n4592 = n4590 & ~n4591;
  assign n4593 = ~n4587 & n4592;
  assign n4594 = n4593 ^ x26;
  assign n4677 = n4676 ^ n4594;
  assign n4584 = n4467 ^ n4400;
  assign n4585 = n4468 & n4584;
  assign n4586 = n4585 ^ n4400;
  assign n4678 = n4677 ^ n4586;
  assign n4576 = n1667 & n1746;
  assign n4577 = x82 & n1871;
  assign n4578 = x83 & n1750;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = x84 & n1873;
  assign n4581 = n4579 & ~n4580;
  assign n4582 = ~n4576 & n4581;
  assign n4583 = n4582 ^ x23;
  assign n4679 = n4678 ^ n4583;
  assign n4573 = n4469 ^ n4389;
  assign n4574 = ~n4470 & ~n4573;
  assign n4575 = n4574 ^ n4389;
  assign n4680 = n4679 ^ n4575;
  assign n4565 = n1404 & n2039;
  assign n4566 = x86 & n1408;
  assign n4567 = x85 & n1514;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = x87 & n1517;
  assign n4570 = n4568 & ~n4569;
  assign n4571 = ~n4565 & n4570;
  assign n4572 = n4571 ^ x20;
  assign n4681 = n4680 ^ n4572;
  assign n4562 = n4471 ^ n4378;
  assign n4563 = n4472 & n4562;
  assign n4564 = n4563 ^ n4378;
  assign n4682 = n4681 ^ n4564;
  assign n4554 = n1098 & n2448;
  assign n4555 = x89 & n1102;
  assign n4556 = x88 & n1198;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = x90 & n1201;
  assign n4559 = n4557 & ~n4558;
  assign n4560 = ~n4554 & n4559;
  assign n4561 = n4560 ^ x17;
  assign n4683 = n4682 ^ n4561;
  assign n4551 = n4473 ^ n4367;
  assign n4552 = ~n4474 & ~n4551;
  assign n4553 = n4552 ^ n4367;
  assign n4684 = n4683 ^ n4553;
  assign n4543 = n821 & n2901;
  assign n4544 = x91 & n898;
  assign n4545 = x93 & n901;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = x92 & n824;
  assign n4548 = n4546 & ~n4547;
  assign n4549 = ~n4543 & n4548;
  assign n4550 = n4549 ^ x14;
  assign n4685 = n4684 ^ n4550;
  assign n4540 = n4475 ^ n4356;
  assign n4541 = n4476 & n4540;
  assign n4542 = n4541 ^ n4356;
  assign n4686 = n4685 ^ n4542;
  assign n4532 = n596 & n3403;
  assign n4533 = x94 & n673;
  assign n4534 = x95 & n601;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = x96 & n676;
  assign n4537 = n4535 & ~n4536;
  assign n4538 = ~n4532 & n4537;
  assign n4539 = n4538 ^ x11;
  assign n4687 = n4686 ^ n4539;
  assign n4529 = n4477 ^ n4345;
  assign n4530 = ~n4478 & ~n4529;
  assign n4531 = n4530 ^ n4345;
  assign n4688 = n4687 ^ n4531;
  assign n4521 = n399 & n3943;
  assign n4522 = x97 & n478;
  assign n4523 = x98 & n402;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = x99 & n470;
  assign n4526 = n4524 & ~n4525;
  assign n4527 = ~n4521 & n4526;
  assign n4528 = n4527 ^ x8;
  assign n4689 = n4688 ^ n4528;
  assign n4518 = n4479 ^ n4334;
  assign n4519 = n4480 & n4518;
  assign n4520 = n4519 ^ n4334;
  assign n4690 = n4689 ^ n4520;
  assign n4509 = n3933 ^ x102;
  assign n4510 = n239 & n4509;
  assign n4511 = x100 & n249;
  assign n4512 = x102 & n280;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = x101 & n242;
  assign n4515 = n4513 & ~n4514;
  assign n4516 = ~n4510 & n4515;
  assign n4517 = n4516 ^ x5;
  assign n4691 = n4690 ^ n4517;
  assign n4506 = n4481 ^ n4322;
  assign n4507 = ~n4482 & n4506;
  assign n4508 = n4507 ^ n4322;
  assign n4692 = n4691 ^ n4508;
  assign n4491 = x104 & ~n4312;
  assign n4492 = ~x104 & ~n4311;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = n169 & ~n4493;
  assign n4495 = n4494 ^ x1;
  assign n4496 = n4495 ^ x105;
  assign n4489 = x1 & x104;
  assign n4490 = n4489 ^ x2;
  assign n4497 = n4496 ^ n4490;
  assign n4498 = n4497 ^ n4496;
  assign n4499 = x103 & n197;
  assign n4500 = n4499 ^ n4496;
  assign n4501 = n4500 ^ n4496;
  assign n4502 = n4498 & ~n4501;
  assign n4503 = n4502 ^ n4496;
  assign n4504 = ~x0 & n4503;
  assign n4505 = n4504 ^ n4496;
  assign n4693 = n4692 ^ n4505;
  assign n4486 = n4483 ^ n4305;
  assign n4487 = n4484 & ~n4486;
  assign n4488 = n4487 ^ n4305;
  assign n4694 = n4693 ^ n4488;
  assign n4859 = ~n4641 & n4659;
  assign n4860 = x41 & ~n4859;
  assign n4850 = x66 & n4646;
  assign n4851 = x65 & n4653;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = n4642 ^ n285;
  assign n4854 = n4853 ^ n285;
  assign n4855 = n2246 & ~n4854;
  assign n4856 = n4855 ^ n285;
  assign n4857 = n4260 & n4856;
  assign n4858 = n4852 & ~n4857;
  assign n4861 = n4860 ^ n4858;
  assign n4848 = x42 ^ x41;
  assign n4849 = x64 & n4848;
  assign n4862 = n4861 ^ n4849;
  assign n4840 = n458 & n4040;
  assign n4841 = x68 & n4267;
  assign n4842 = x69 & n4044;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = x70 & n4270;
  assign n4845 = n4843 & ~n4844;
  assign n4846 = ~n4840 & n4845;
  assign n4847 = n4846 ^ x38;
  assign n4863 = n4862 ^ n4847;
  assign n4837 = n4668 ^ n4630;
  assign n4838 = ~n4669 & ~n4837;
  assign n4839 = n4838 ^ n4630;
  assign n4864 = n4863 ^ n4839;
  assign n4829 = ~n653 & n3522;
  assign n4830 = x72 & n3526;
  assign n4831 = x71 & n3699;
  assign n4832 = ~n4830 & ~n4831;
  assign n4833 = x73 & n3701;
  assign n4834 = n4832 & ~n4833;
  assign n4835 = ~n4829 & n4834;
  assign n4836 = n4835 ^ x35;
  assign n4865 = n4864 ^ n4836;
  assign n4826 = n4670 ^ n4619;
  assign n4827 = n4671 & n4826;
  assign n4828 = n4827 ^ n4619;
  assign n4866 = n4865 ^ n4828;
  assign n4818 = n870 & n3009;
  assign n4819 = x74 & n3181;
  assign n4820 = x75 & n3013;
  assign n4821 = ~n4819 & ~n4820;
  assign n4822 = x76 & n3183;
  assign n4823 = n4821 & ~n4822;
  assign n4824 = ~n4818 & n4823;
  assign n4825 = n4824 ^ x32;
  assign n4867 = n4866 ^ n4825;
  assign n4815 = n4672 ^ n4608;
  assign n4816 = ~n4673 & ~n4815;
  assign n4817 = n4816 ^ n4608;
  assign n4868 = n4867 ^ n4817;
  assign n4807 = n1149 & n2527;
  assign n4808 = x77 & n2690;
  assign n4809 = x79 & n2693;
  assign n4810 = ~n4808 & ~n4809;
  assign n4811 = x78 & n2530;
  assign n4812 = n4810 & ~n4811;
  assign n4813 = ~n4807 & n4812;
  assign n4814 = n4813 ^ x29;
  assign n4869 = n4868 ^ n4814;
  assign n4804 = n4674 ^ n4597;
  assign n4805 = n4675 & n4804;
  assign n4806 = n4805 ^ n4597;
  assign n4870 = n4869 ^ n4806;
  assign n4796 = n1454 & n2102;
  assign n4797 = x81 & n2105;
  assign n4798 = x80 & n2112;
  assign n4799 = ~n4797 & ~n4798;
  assign n4800 = x82 & n2381;
  assign n4801 = n4799 & ~n4800;
  assign n4802 = ~n4796 & n4801;
  assign n4803 = n4802 ^ x26;
  assign n4871 = n4870 ^ n4803;
  assign n4793 = n4676 ^ n4586;
  assign n4794 = ~n4677 & ~n4793;
  assign n4795 = n4794 ^ n4586;
  assign n4872 = n4871 ^ n4795;
  assign n4785 = n1746 & n1801;
  assign n4786 = x83 & n1871;
  assign n4787 = x84 & n1750;
  assign n4788 = ~n4786 & ~n4787;
  assign n4789 = x85 & n1873;
  assign n4790 = n4788 & ~n4789;
  assign n4791 = ~n4785 & n4790;
  assign n4792 = n4791 ^ x23;
  assign n4873 = n4872 ^ n4792;
  assign n4782 = n4678 ^ n4575;
  assign n4783 = n4679 & n4782;
  assign n4784 = n4783 ^ n4575;
  assign n4874 = n4873 ^ n4784;
  assign n4774 = n1404 & n2176;
  assign n4775 = x87 & n1408;
  assign n4776 = x86 & n1514;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = x88 & n1517;
  assign n4779 = n4777 & ~n4778;
  assign n4780 = ~n4774 & n4779;
  assign n4781 = n4780 ^ x20;
  assign n4875 = n4874 ^ n4781;
  assign n4771 = n4680 ^ n4564;
  assign n4772 = ~n4681 & ~n4771;
  assign n4773 = n4772 ^ n4564;
  assign n4876 = n4875 ^ n4773;
  assign n4763 = n1098 & n2607;
  assign n4764 = x90 & n1102;
  assign n4765 = x89 & n1198;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = x91 & n1201;
  assign n4768 = n4766 & ~n4767;
  assign n4769 = ~n4763 & n4768;
  assign n4770 = n4769 ^ x17;
  assign n4877 = n4876 ^ n4770;
  assign n4760 = n4682 ^ n4553;
  assign n4761 = n4683 & n4760;
  assign n4762 = n4761 ^ n4553;
  assign n4878 = n4877 ^ n4762;
  assign n4752 = n821 & n3078;
  assign n4753 = x92 & n898;
  assign n4754 = x93 & n824;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = x94 & n901;
  assign n4757 = n4755 & ~n4756;
  assign n4758 = ~n4752 & n4757;
  assign n4759 = n4758 ^ x14;
  assign n4879 = n4878 ^ n4759;
  assign n4749 = n4684 ^ n4542;
  assign n4750 = ~n4685 & ~n4749;
  assign n4751 = n4750 ^ n4542;
  assign n4880 = n4879 ^ n4751;
  assign n4741 = n596 & n3585;
  assign n4742 = x95 & n673;
  assign n4743 = x96 & n601;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = x97 & n676;
  assign n4746 = n4744 & ~n4745;
  assign n4747 = ~n4741 & n4746;
  assign n4748 = n4747 ^ x11;
  assign n4881 = n4880 ^ n4748;
  assign n4738 = n4686 ^ n4531;
  assign n4739 = n4687 & n4738;
  assign n4740 = n4739 ^ n4531;
  assign n4882 = n4881 ^ n4740;
  assign n4730 = n399 & n4141;
  assign n4731 = x98 & n478;
  assign n4732 = x100 & n470;
  assign n4733 = ~n4731 & ~n4732;
  assign n4734 = x99 & n402;
  assign n4735 = n4733 & ~n4734;
  assign n4736 = ~n4730 & n4735;
  assign n4737 = n4736 ^ x8;
  assign n4883 = n4882 ^ n4737;
  assign n4727 = n4688 ^ n4520;
  assign n4728 = ~n4689 & ~n4727;
  assign n4729 = n4728 ^ n4520;
  assign n4884 = n4883 ^ n4729;
  assign n4718 = n4131 ^ x103;
  assign n4719 = n239 & n4718;
  assign n4720 = x101 & n249;
  assign n4721 = x103 & n280;
  assign n4722 = ~n4720 & ~n4721;
  assign n4723 = x102 & n242;
  assign n4724 = n4722 & ~n4723;
  assign n4725 = ~n4719 & n4724;
  assign n4726 = n4725 ^ x5;
  assign n4885 = n4884 ^ n4726;
  assign n4715 = n4690 ^ n4508;
  assign n4716 = n4691 & ~n4715;
  assign n4717 = n4716 ^ n4508;
  assign n4886 = n4885 ^ n4717;
  assign n4704 = x105 ^ x2;
  assign n4705 = n4704 ^ x104;
  assign n4706 = n4705 ^ n4704;
  assign n4707 = n4704 ^ x105;
  assign n4708 = ~n4706 & n4707;
  assign n4709 = n4708 ^ n4704;
  assign n4710 = ~x1 & n4709;
  assign n4711 = n4710 ^ n4704;
  assign n4698 = x105 & ~n4492;
  assign n4699 = ~x105 & ~n4491;
  assign n4700 = ~n4698 & ~n4699;
  assign n4701 = n169 & ~n4700;
  assign n4702 = n4701 ^ x1;
  assign n4703 = n4702 ^ x106;
  assign n4712 = n4711 ^ n4703;
  assign n4713 = ~x0 & n4712;
  assign n4714 = n4713 ^ n4703;
  assign n4887 = n4886 ^ n4714;
  assign n4695 = n4692 ^ n4488;
  assign n4696 = ~n4693 & n4695;
  assign n4697 = n4696 ^ n4488;
  assign n4888 = n4887 ^ n4697;
  assign n5059 = ~n4849 & ~n4861;
  assign n5060 = n4858 ^ x41;
  assign n5061 = ~n5059 & ~n5060;
  assign n5054 = x65 ^ x42;
  assign n5055 = n4848 & ~n5054;
  assign n5056 = n5055 ^ x41;
  assign n5057 = n5056 ^ x43;
  assign n5051 = x41 & x42;
  assign n5052 = n5051 ^ x43;
  assign n5053 = ~x64 & n5052;
  assign n5058 = n5057 ^ n5053;
  assign n5062 = n5061 ^ n5058;
  assign n5042 = n321 & n4643;
  assign n5043 = x67 & n4646;
  assign n5044 = x66 & n4653;
  assign n5045 = ~n5043 & ~n5044;
  assign n5046 = n4260 & ~n4642;
  assign n5047 = x68 & n5046;
  assign n5048 = n5045 & ~n5047;
  assign n5049 = ~n5042 & n5048;
  assign n5050 = n5049 ^ x41;
  assign n5063 = n5062 ^ n5050;
  assign n5034 = n517 & n4040;
  assign n5035 = x69 & n4267;
  assign n5036 = x70 & n4044;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = x71 & n4270;
  assign n5039 = n5037 & ~n5038;
  assign n5040 = ~n5034 & n5039;
  assign n5041 = n5040 ^ x38;
  assign n5064 = n5063 ^ n5041;
  assign n5031 = n4862 ^ n4839;
  assign n5032 = ~n4863 & ~n5031;
  assign n5033 = n5032 ^ n4839;
  assign n5065 = n5064 ^ n5033;
  assign n5023 = ~n721 & n3522;
  assign n5024 = x73 & n3526;
  assign n5025 = x72 & n3699;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = x74 & n3701;
  assign n5028 = n5026 & ~n5027;
  assign n5029 = ~n5023 & n5028;
  assign n5030 = n5029 ^ x35;
  assign n5066 = n5065 ^ n5030;
  assign n5020 = n4864 ^ n4828;
  assign n5021 = n4865 & n5020;
  assign n5022 = n5021 ^ n4828;
  assign n5067 = n5066 ^ n5022;
  assign n5012 = n956 & n3009;
  assign n5013 = x75 & n3181;
  assign n5014 = x76 & n3013;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = x77 & n3183;
  assign n5017 = n5015 & ~n5016;
  assign n5018 = ~n5012 & n5017;
  assign n5019 = n5018 ^ x32;
  assign n5068 = n5067 ^ n5019;
  assign n5009 = n4866 ^ n4817;
  assign n5010 = ~n4867 & ~n5009;
  assign n5011 = n5010 ^ n4817;
  assign n5069 = n5068 ^ n5011;
  assign n5001 = n1242 & n2527;
  assign n5002 = x78 & n2690;
  assign n5003 = x79 & n2530;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = x80 & n2693;
  assign n5006 = n5004 & ~n5005;
  assign n5007 = ~n5001 & n5006;
  assign n5008 = n5007 ^ x29;
  assign n5070 = n5069 ^ n5008;
  assign n4998 = n4868 ^ n4806;
  assign n4999 = n4869 & n4998;
  assign n5000 = n4999 ^ n4806;
  assign n5071 = n5070 ^ n5000;
  assign n4990 = n1560 & n2102;
  assign n4991 = x81 & n2112;
  assign n4992 = x82 & n2105;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = x83 & n2381;
  assign n4995 = n4993 & ~n4994;
  assign n4996 = ~n4990 & n4995;
  assign n4997 = n4996 ^ x26;
  assign n5072 = n5071 ^ n4997;
  assign n4987 = n4870 ^ n4795;
  assign n4988 = ~n4871 & ~n4987;
  assign n4989 = n4988 ^ n4795;
  assign n5073 = n5072 ^ n4989;
  assign n4979 = n1746 & n1920;
  assign n4980 = x84 & n1871;
  assign n4981 = x85 & n1750;
  assign n4982 = ~n4980 & ~n4981;
  assign n4983 = x86 & n1873;
  assign n4984 = n4982 & ~n4983;
  assign n4985 = ~n4979 & n4984;
  assign n4986 = n4985 ^ x23;
  assign n5074 = n5073 ^ n4986;
  assign n4976 = n4872 ^ n4784;
  assign n4977 = n4873 & n4976;
  assign n4978 = n4977 ^ n4784;
  assign n5075 = n5074 ^ n4978;
  assign n4968 = n1404 & n2310;
  assign n4969 = x87 & n1514;
  assign n4970 = x88 & n1408;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = x89 & n1517;
  assign n4973 = n4971 & ~n4972;
  assign n4974 = ~n4968 & n4973;
  assign n4975 = n4974 ^ x20;
  assign n5076 = n5075 ^ n4975;
  assign n4965 = n4874 ^ n4773;
  assign n4966 = ~n4875 & ~n4965;
  assign n4967 = n4966 ^ n4773;
  assign n5077 = n5076 ^ n4967;
  assign n4957 = n1098 & n2755;
  assign n4958 = x90 & n1198;
  assign n4959 = x91 & n1102;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = x92 & n1201;
  assign n4962 = n4960 & ~n4961;
  assign n4963 = ~n4957 & n4962;
  assign n4964 = n4963 ^ x17;
  assign n5078 = n5077 ^ n4964;
  assign n4954 = n4876 ^ n4762;
  assign n4955 = n4877 & n4954;
  assign n4956 = n4955 ^ n4762;
  assign n5079 = n5078 ^ n4956;
  assign n4946 = n821 & n3247;
  assign n4947 = x93 & n898;
  assign n4948 = x94 & n824;
  assign n4949 = ~n4947 & ~n4948;
  assign n4950 = x95 & n901;
  assign n4951 = n4949 & ~n4950;
  assign n4952 = ~n4946 & n4951;
  assign n4953 = n4952 ^ x14;
  assign n5080 = n5079 ^ n4953;
  assign n4943 = n4878 ^ n4751;
  assign n4944 = ~n4879 & ~n4943;
  assign n4945 = n4944 ^ n4751;
  assign n5081 = n5080 ^ n4945;
  assign n4935 = n596 & n3763;
  assign n4936 = x97 & n601;
  assign n4937 = x98 & n676;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = x96 & n673;
  assign n4940 = n4938 & ~n4939;
  assign n4941 = ~n4935 & n4940;
  assign n4942 = n4941 ^ x11;
  assign n5082 = n5081 ^ n4942;
  assign n4932 = n4880 ^ n4740;
  assign n4933 = n4881 & n4932;
  assign n4934 = n4933 ^ n4740;
  assign n5083 = n5082 ^ n4934;
  assign n4924 = n399 & n4323;
  assign n4925 = x99 & n478;
  assign n4926 = x100 & n402;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = x101 & n470;
  assign n4929 = n4927 & ~n4928;
  assign n4930 = ~n4924 & n4929;
  assign n4931 = n4930 ^ x8;
  assign n5084 = n5083 ^ n4931;
  assign n4921 = n4882 ^ n4729;
  assign n4922 = ~n4883 & ~n4921;
  assign n4923 = n4922 ^ n4729;
  assign n5085 = n5084 ^ n4923;
  assign n4912 = n4313 ^ x104;
  assign n4913 = n239 & n4912;
  assign n4914 = x102 & n249;
  assign n4915 = x103 & n242;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = x104 & n280;
  assign n4918 = n4916 & ~n4917;
  assign n4919 = ~n4913 & n4918;
  assign n4920 = n4919 ^ x5;
  assign n5086 = n5085 ^ n4920;
  assign n4909 = n4884 ^ n4717;
  assign n4910 = n4885 & ~n4909;
  assign n4911 = n4910 ^ n4717;
  assign n5087 = n5086 ^ n4911;
  assign n4894 = ~x106 & ~n4698;
  assign n4895 = x106 & ~n4699;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = n169 & ~n4896;
  assign n4898 = n4897 ^ x1;
  assign n4899 = n4898 ^ x107;
  assign n4892 = x106 ^ x2;
  assign n4893 = x1 & n4892;
  assign n4900 = n4899 ^ n4893;
  assign n4901 = n4900 ^ n4899;
  assign n4902 = ~x105 & n197;
  assign n4903 = n4902 ^ n4899;
  assign n4904 = n4903 ^ n4899;
  assign n4905 = ~n4901 & ~n4904;
  assign n4906 = n4905 ^ n4899;
  assign n4907 = ~x0 & ~n4906;
  assign n4908 = n4907 ^ n4899;
  assign n5088 = n5087 ^ n4908;
  assign n4889 = n4886 ^ n4697;
  assign n4890 = ~n4887 & n4889;
  assign n4891 = n4890 ^ n4697;
  assign n5089 = n5088 ^ n4891;
  assign n5288 = n789 & n3522;
  assign n5289 = x73 & n3699;
  assign n5290 = x75 & n3701;
  assign n5291 = ~n5289 & ~n5290;
  assign n5292 = x74 & n3526;
  assign n5293 = n5291 & ~n5292;
  assign n5294 = ~n5288 & n5293;
  assign n5295 = n5294 ^ x35;
  assign n5285 = n5065 ^ n5022;
  assign n5286 = n5066 & n5285;
  assign n5287 = n5286 ^ n5022;
  assign n5296 = n5295 ^ n5287;
  assign n5247 = ~x41 & ~x42;
  assign n5258 = ~x43 & x44;
  assign n5259 = n5247 & n5258;
  assign n5260 = x64 & n5259;
  assign n5261 = x44 ^ x43;
  assign n5262 = n4848 & n5261;
  assign n5263 = n142 & n5262;
  assign n5264 = n5247 ^ n5051;
  assign n5265 = x43 & n5264;
  assign n5266 = n5265 ^ n5051;
  assign n5267 = ~n5263 & ~n5266;
  assign n5268 = x65 & ~n5267;
  assign n5269 = n152 & n5261;
  assign n5270 = x66 & n4848;
  assign n5271 = ~n5269 & n5270;
  assign n5272 = ~n5268 & ~n5271;
  assign n5273 = n5272 ^ x44;
  assign n5274 = x43 & x64;
  assign n5275 = n5051 & n5274;
  assign n5276 = n5272 & n5275;
  assign n5277 = n5273 & n5276;
  assign n5278 = n5277 ^ n5273;
  assign n5279 = ~n5260 & ~n5278;
  assign n5248 = ~n233 & ~n5247;
  assign n5249 = n5248 ^ n5051;
  assign n5250 = x64 ^ x43;
  assign n5251 = n5250 ^ x43;
  assign n5252 = n5248 ^ x43;
  assign n5253 = ~n5251 & n5252;
  assign n5254 = n5253 ^ x43;
  assign n5255 = ~n5249 & ~n5254;
  assign n5256 = n5255 ^ n5051;
  assign n5257 = x44 & n5256;
  assign n5280 = n5279 ^ n5257;
  assign n5239 = n420 & n4643;
  assign n5240 = x67 & n4653;
  assign n5241 = x68 & n4646;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = x69 & n5046;
  assign n5244 = n5242 & ~n5243;
  assign n5245 = ~n5239 & n5244;
  assign n5246 = n5245 ^ x41;
  assign n5281 = n5280 ^ n5246;
  assign n5236 = n5058 ^ n5050;
  assign n5237 = n5062 & n5236;
  assign n5238 = n5237 ^ n5061;
  assign n5282 = n5281 ^ n5238;
  assign n5228 = n575 & n4040;
  assign n5229 = x71 & n4044;
  assign n5230 = x70 & n4267;
  assign n5231 = ~n5229 & ~n5230;
  assign n5232 = x72 & n4270;
  assign n5233 = n5231 & ~n5232;
  assign n5234 = ~n5228 & n5233;
  assign n5235 = n5234 ^ x38;
  assign n5283 = n5282 ^ n5235;
  assign n5225 = n5063 ^ n5033;
  assign n5226 = ~n5064 & ~n5225;
  assign n5227 = n5226 ^ n5033;
  assign n5284 = n5283 ^ n5227;
  assign n5297 = n5296 ^ n5284;
  assign n5217 = n1041 & n3009;
  assign n5218 = x76 & n3181;
  assign n5219 = x77 & n3013;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = x78 & n3183;
  assign n5222 = n5220 & ~n5221;
  assign n5223 = ~n5217 & n5222;
  assign n5224 = n5223 ^ x32;
  assign n5298 = n5297 ^ n5224;
  assign n5214 = n5067 ^ n5011;
  assign n5215 = ~n5068 & ~n5214;
  assign n5216 = n5215 ^ n5011;
  assign n5299 = n5298 ^ n5216;
  assign n5206 = n1340 & n2527;
  assign n5207 = x79 & n2690;
  assign n5208 = x80 & n2530;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = x81 & n2693;
  assign n5211 = n5209 & ~n5210;
  assign n5212 = ~n5206 & n5211;
  assign n5213 = n5212 ^ x29;
  assign n5300 = n5299 ^ n5213;
  assign n5203 = n5069 ^ n5000;
  assign n5204 = n5070 & n5203;
  assign n5205 = n5204 ^ n5000;
  assign n5301 = n5300 ^ n5205;
  assign n5195 = n1667 & n2102;
  assign n5196 = x82 & n2112;
  assign n5197 = x84 & n2381;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = x83 & n2105;
  assign n5200 = n5198 & ~n5199;
  assign n5201 = ~n5195 & n5200;
  assign n5202 = n5201 ^ x26;
  assign n5302 = n5301 ^ n5202;
  assign n5192 = n5071 ^ n4989;
  assign n5193 = ~n5072 & ~n5192;
  assign n5194 = n5193 ^ n4989;
  assign n5303 = n5302 ^ n5194;
  assign n5184 = n1746 & n2039;
  assign n5185 = x85 & n1871;
  assign n5186 = x86 & n1750;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = x87 & n1873;
  assign n5189 = n5187 & ~n5188;
  assign n5190 = ~n5184 & n5189;
  assign n5191 = n5190 ^ x23;
  assign n5304 = n5303 ^ n5191;
  assign n5181 = n5073 ^ n4978;
  assign n5182 = n5074 & n5181;
  assign n5183 = n5182 ^ n4978;
  assign n5305 = n5304 ^ n5183;
  assign n5173 = n1404 & n2448;
  assign n5174 = x89 & n1408;
  assign n5175 = x88 & n1514;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = x90 & n1517;
  assign n5178 = n5176 & ~n5177;
  assign n5179 = ~n5173 & n5178;
  assign n5180 = n5179 ^ x20;
  assign n5306 = n5305 ^ n5180;
  assign n5170 = n5075 ^ n4967;
  assign n5171 = ~n5076 & ~n5170;
  assign n5172 = n5171 ^ n4967;
  assign n5307 = n5306 ^ n5172;
  assign n5162 = n1098 & n2901;
  assign n5163 = x92 & n1102;
  assign n5164 = x91 & n1198;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = x93 & n1201;
  assign n5167 = n5165 & ~n5166;
  assign n5168 = ~n5162 & n5167;
  assign n5169 = n5168 ^ x17;
  assign n5308 = n5307 ^ n5169;
  assign n5159 = n5077 ^ n4956;
  assign n5160 = n5078 & n5159;
  assign n5161 = n5160 ^ n4956;
  assign n5309 = n5308 ^ n5161;
  assign n5151 = n821 & n3403;
  assign n5152 = x94 & n898;
  assign n5153 = x96 & n901;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = x95 & n824;
  assign n5156 = n5154 & ~n5155;
  assign n5157 = ~n5151 & n5156;
  assign n5158 = n5157 ^ x14;
  assign n5310 = n5309 ^ n5158;
  assign n5148 = n5079 ^ n4945;
  assign n5149 = ~n5080 & ~n5148;
  assign n5150 = n5149 ^ n4945;
  assign n5311 = n5310 ^ n5150;
  assign n5140 = n596 & n3943;
  assign n5141 = x97 & n673;
  assign n5142 = x99 & n676;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = x98 & n601;
  assign n5145 = n5143 & ~n5144;
  assign n5146 = ~n5140 & n5145;
  assign n5147 = n5146 ^ x11;
  assign n5312 = n5311 ^ n5147;
  assign n5137 = n5081 ^ n4934;
  assign n5138 = n5082 & n5137;
  assign n5139 = n5138 ^ n4934;
  assign n5313 = n5312 ^ n5139;
  assign n5129 = n399 & n4509;
  assign n5130 = x100 & n478;
  assign n5131 = x101 & n402;
  assign n5132 = ~n5130 & ~n5131;
  assign n5133 = x102 & n470;
  assign n5134 = n5132 & ~n5133;
  assign n5135 = ~n5129 & n5134;
  assign n5136 = n5135 ^ x8;
  assign n5314 = n5313 ^ n5136;
  assign n5126 = n5083 ^ n4923;
  assign n5127 = ~n5084 & ~n5126;
  assign n5128 = n5127 ^ n4923;
  assign n5315 = n5314 ^ n5128;
  assign n5117 = n4493 ^ x105;
  assign n5118 = n239 & n5117;
  assign n5119 = x103 & n249;
  assign n5120 = x104 & n242;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = x105 & n280;
  assign n5123 = n5121 & ~n5122;
  assign n5124 = ~n5118 & n5123;
  assign n5125 = n5124 ^ x5;
  assign n5316 = n5315 ^ n5125;
  assign n5114 = n5085 ^ n4911;
  assign n5115 = n5086 & ~n5114;
  assign n5116 = n5115 ^ n4911;
  assign n5317 = n5316 ^ n5116;
  assign n5101 = x107 ^ x106;
  assign n5102 = n4699 ^ n4698;
  assign n5103 = n4698 ^ x107;
  assign n5104 = n5103 ^ n4698;
  assign n5105 = n5102 & ~n5104;
  assign n5106 = n5105 ^ n4698;
  assign n5107 = n5101 & ~n5106;
  assign n5108 = n169 & ~n5107;
  assign n5109 = n5108 ^ x1;
  assign n5110 = n5109 ^ x108;
  assign n5093 = x107 ^ x2;
  assign n5094 = n5093 ^ x106;
  assign n5095 = n5094 ^ n5093;
  assign n5096 = n5093 ^ x107;
  assign n5097 = ~n5095 & n5096;
  assign n5098 = n5097 ^ n5093;
  assign n5099 = ~x1 & n5098;
  assign n5100 = n5099 ^ n5093;
  assign n5111 = n5110 ^ n5100;
  assign n5112 = ~x0 & n5111;
  assign n5113 = n5112 ^ n5110;
  assign n5318 = n5317 ^ n5113;
  assign n5090 = n5087 ^ n4891;
  assign n5091 = ~n5088 & n5090;
  assign n5092 = n5091 ^ n4891;
  assign n5319 = n5318 ^ n5092;
  assign n5505 = ~n653 & n4040;
  assign n5506 = x71 & n4267;
  assign n5507 = x73 & n4270;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = x72 & n4044;
  assign n5510 = n5508 & ~n5509;
  assign n5511 = ~n5505 & n5510;
  assign n5512 = n5511 ^ x38;
  assign n5502 = n5282 ^ n5227;
  assign n5503 = ~n5283 & ~n5502;
  assign n5504 = n5503 ^ n5227;
  assign n5513 = n5512 ^ n5504;
  assign n5498 = n5257 & n5279;
  assign n5483 = x66 & n5266;
  assign n5484 = n5051 ^ x44;
  assign n5485 = n5484 ^ n5051;
  assign n5486 = n5264 & n5485;
  assign n5487 = n5486 ^ n5051;
  assign n5488 = n5261 & n5487;
  assign n5489 = x65 & n5488;
  assign n5490 = ~n5483 & ~n5489;
  assign n5491 = n4848 & ~n5261;
  assign n5492 = x67 & n5491;
  assign n5493 = n5490 & ~n5492;
  assign n5494 = n285 & n5262;
  assign n5495 = n5493 & ~n5494;
  assign n5496 = n5495 ^ x44;
  assign n5481 = x45 ^ x44;
  assign n5482 = x64 & n5481;
  assign n5497 = n5496 ^ n5482;
  assign n5499 = n5498 ^ n5497;
  assign n5473 = n458 & n4643;
  assign n5474 = x69 & n4646;
  assign n5475 = x68 & n4653;
  assign n5476 = ~n5474 & ~n5475;
  assign n5477 = x70 & n5046;
  assign n5478 = n5476 & ~n5477;
  assign n5479 = ~n5473 & n5478;
  assign n5480 = n5479 ^ x41;
  assign n5500 = n5499 ^ n5480;
  assign n5470 = n5280 ^ n5238;
  assign n5471 = n5281 & n5470;
  assign n5472 = n5471 ^ n5238;
  assign n5501 = n5500 ^ n5472;
  assign n5514 = n5513 ^ n5501;
  assign n5462 = n870 & n3522;
  assign n5463 = x74 & n3699;
  assign n5464 = x76 & n3701;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = x75 & n3526;
  assign n5467 = n5465 & ~n5466;
  assign n5468 = ~n5462 & n5467;
  assign n5469 = n5468 ^ x35;
  assign n5515 = n5514 ^ n5469;
  assign n5459 = n5295 ^ n5284;
  assign n5460 = ~n5296 & n5459;
  assign n5461 = n5460 ^ n5287;
  assign n5516 = n5515 ^ n5461;
  assign n5451 = n1149 & n3009;
  assign n5452 = x77 & n3181;
  assign n5453 = x78 & n3013;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = x79 & n3183;
  assign n5456 = n5454 & ~n5455;
  assign n5457 = ~n5451 & n5456;
  assign n5458 = n5457 ^ x32;
  assign n5517 = n5516 ^ n5458;
  assign n5448 = n5297 ^ n5216;
  assign n5449 = ~n5298 & ~n5448;
  assign n5450 = n5449 ^ n5216;
  assign n5518 = n5517 ^ n5450;
  assign n5440 = n1454 & n2527;
  assign n5441 = x80 & n2690;
  assign n5442 = x81 & n2530;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = x82 & n2693;
  assign n5445 = n5443 & ~n5444;
  assign n5446 = ~n5440 & n5445;
  assign n5447 = n5446 ^ x29;
  assign n5519 = n5518 ^ n5447;
  assign n5437 = n5299 ^ n5205;
  assign n5438 = n5300 & n5437;
  assign n5439 = n5438 ^ n5205;
  assign n5520 = n5519 ^ n5439;
  assign n5429 = n1801 & n2102;
  assign n5430 = x83 & n2112;
  assign n5431 = x85 & n2381;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = x84 & n2105;
  assign n5434 = n5432 & ~n5433;
  assign n5435 = ~n5429 & n5434;
  assign n5436 = n5435 ^ x26;
  assign n5521 = n5520 ^ n5436;
  assign n5426 = n5301 ^ n5194;
  assign n5427 = ~n5302 & ~n5426;
  assign n5428 = n5427 ^ n5194;
  assign n5522 = n5521 ^ n5428;
  assign n5418 = n1746 & n2176;
  assign n5419 = x86 & n1871;
  assign n5420 = x87 & n1750;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = x88 & n1873;
  assign n5423 = n5421 & ~n5422;
  assign n5424 = ~n5418 & n5423;
  assign n5425 = n5424 ^ x23;
  assign n5523 = n5522 ^ n5425;
  assign n5415 = n5303 ^ n5183;
  assign n5416 = n5304 & n5415;
  assign n5417 = n5416 ^ n5183;
  assign n5524 = n5523 ^ n5417;
  assign n5407 = n1404 & n2607;
  assign n5408 = x89 & n1514;
  assign n5409 = x91 & n1517;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = x90 & n1408;
  assign n5412 = n5410 & ~n5411;
  assign n5413 = ~n5407 & n5412;
  assign n5414 = n5413 ^ x20;
  assign n5525 = n5524 ^ n5414;
  assign n5404 = n5305 ^ n5172;
  assign n5405 = ~n5306 & ~n5404;
  assign n5406 = n5405 ^ n5172;
  assign n5526 = n5525 ^ n5406;
  assign n5396 = n1098 & n3078;
  assign n5397 = x93 & n1102;
  assign n5398 = x92 & n1198;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = x94 & n1201;
  assign n5401 = n5399 & ~n5400;
  assign n5402 = ~n5396 & n5401;
  assign n5403 = n5402 ^ x17;
  assign n5527 = n5526 ^ n5403;
  assign n5393 = n5307 ^ n5161;
  assign n5394 = n5308 & n5393;
  assign n5395 = n5394 ^ n5161;
  assign n5528 = n5527 ^ n5395;
  assign n5385 = n821 & n3585;
  assign n5386 = x95 & n898;
  assign n5387 = x97 & n901;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = x96 & n824;
  assign n5390 = n5388 & ~n5389;
  assign n5391 = ~n5385 & n5390;
  assign n5392 = n5391 ^ x14;
  assign n5529 = n5528 ^ n5392;
  assign n5382 = n5309 ^ n5150;
  assign n5383 = ~n5310 & ~n5382;
  assign n5384 = n5383 ^ n5150;
  assign n5530 = n5529 ^ n5384;
  assign n5374 = n596 & n4141;
  assign n5375 = x98 & n673;
  assign n5376 = x100 & n676;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = x99 & n601;
  assign n5379 = n5377 & ~n5378;
  assign n5380 = ~n5374 & n5379;
  assign n5381 = n5380 ^ x11;
  assign n5531 = n5530 ^ n5381;
  assign n5371 = n5311 ^ n5139;
  assign n5372 = n5312 & n5371;
  assign n5373 = n5372 ^ n5139;
  assign n5532 = n5531 ^ n5373;
  assign n5363 = n399 & n4718;
  assign n5364 = x101 & n478;
  assign n5365 = x102 & n402;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = x103 & n470;
  assign n5368 = n5366 & ~n5367;
  assign n5369 = ~n5363 & n5368;
  assign n5370 = n5369 ^ x8;
  assign n5533 = n5532 ^ n5370;
  assign n5360 = n5313 ^ n5128;
  assign n5361 = ~n5314 & ~n5360;
  assign n5362 = n5361 ^ n5128;
  assign n5534 = n5533 ^ n5362;
  assign n5351 = n4700 ^ x106;
  assign n5352 = n239 & n5351;
  assign n5353 = x104 & n249;
  assign n5354 = x105 & n242;
  assign n5355 = ~n5353 & ~n5354;
  assign n5356 = x106 & n280;
  assign n5357 = n5355 & ~n5356;
  assign n5358 = ~n5352 & n5357;
  assign n5359 = n5358 ^ x5;
  assign n5535 = n5534 ^ n5359;
  assign n5348 = n5315 ^ n5116;
  assign n5349 = n5316 & ~n5348;
  assign n5350 = n5349 ^ n5116;
  assign n5536 = n5535 ^ n5350;
  assign n5335 = x108 ^ x107;
  assign n5336 = n4895 ^ n4894;
  assign n5337 = n4894 ^ x108;
  assign n5338 = n5337 ^ n4894;
  assign n5339 = n5336 & n5338;
  assign n5340 = n5339 ^ n4894;
  assign n5341 = n5335 & ~n5340;
  assign n5342 = n169 & ~n5341;
  assign n5343 = n5342 ^ x1;
  assign n5344 = n5343 ^ x109;
  assign n5323 = x108 ^ x2;
  assign n5324 = n5323 ^ x1;
  assign n5325 = n5324 ^ n5323;
  assign n5326 = n5325 ^ x0;
  assign n5327 = n5323 ^ x108;
  assign n5328 = n5327 ^ x107;
  assign n5329 = ~x107 & ~n5328;
  assign n5330 = n5329 ^ n5323;
  assign n5331 = n5330 ^ x107;
  assign n5332 = n5326 & ~n5331;
  assign n5333 = n5332 ^ n5329;
  assign n5334 = n5333 ^ x107;
  assign n5345 = n5344 ^ n5334;
  assign n5346 = ~x0 & ~n5345;
  assign n5347 = n5346 ^ n5344;
  assign n5537 = n5536 ^ n5347;
  assign n5320 = n5317 ^ n5092;
  assign n5321 = ~n5318 & n5320;
  assign n5322 = n5321 ^ n5092;
  assign n5538 = n5537 ^ n5322;
  assign n5735 = n956 & n3522;
  assign n5736 = x75 & n3699;
  assign n5737 = x76 & n3526;
  assign n5738 = ~n5736 & ~n5737;
  assign n5739 = x77 & n3701;
  assign n5740 = n5738 & ~n5739;
  assign n5741 = ~n5735 & n5740;
  assign n5742 = n5741 ^ x35;
  assign n5732 = n5514 ^ n5461;
  assign n5733 = ~n5515 & ~n5732;
  assign n5734 = n5733 ^ n5461;
  assign n5743 = n5742 ^ n5734;
  assign n5720 = n517 & n4643;
  assign n5721 = x70 & n4646;
  assign n5722 = x69 & n4653;
  assign n5723 = ~n5721 & ~n5722;
  assign n5724 = x71 & n5046;
  assign n5725 = n5723 & ~n5724;
  assign n5726 = ~n5720 & n5725;
  assign n5727 = n5726 ^ x41;
  assign n5717 = n5499 ^ n5472;
  assign n5718 = ~n5500 & ~n5717;
  assign n5719 = n5718 ^ n5472;
  assign n5728 = n5727 ^ n5719;
  assign n5714 = ~n5482 & ~n5498;
  assign n5715 = ~n5496 & ~n5714;
  assign n5709 = x44 & x45;
  assign n5710 = n5709 ^ x46;
  assign n5711 = ~x64 & n5710;
  assign n5705 = x65 ^ x45;
  assign n5706 = n5481 & ~n5705;
  assign n5707 = n5706 ^ x44;
  assign n5708 = n5707 ^ x46;
  assign n5712 = n5711 ^ n5708;
  assign n5697 = n321 & n5262;
  assign n5698 = x67 & n5266;
  assign n5699 = x66 & n5488;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = x68 & n5491;
  assign n5702 = n5700 & ~n5701;
  assign n5703 = ~n5697 & n5702;
  assign n5704 = n5703 ^ x44;
  assign n5713 = n5712 ^ n5704;
  assign n5716 = n5715 ^ n5713;
  assign n5729 = n5728 ^ n5716;
  assign n5689 = ~n721 & n4040;
  assign n5690 = x73 & n4044;
  assign n5691 = x72 & n4267;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = x74 & n4270;
  assign n5694 = n5692 & ~n5693;
  assign n5695 = ~n5689 & n5694;
  assign n5696 = n5695 ^ x38;
  assign n5730 = n5729 ^ n5696;
  assign n5686 = n5512 ^ n5501;
  assign n5687 = ~n5513 & n5686;
  assign n5688 = n5687 ^ n5504;
  assign n5731 = n5730 ^ n5688;
  assign n5744 = n5743 ^ n5731;
  assign n5678 = n1242 & n3009;
  assign n5679 = x79 & n3013;
  assign n5680 = x78 & n3181;
  assign n5681 = ~n5679 & ~n5680;
  assign n5682 = x80 & n3183;
  assign n5683 = n5681 & ~n5682;
  assign n5684 = ~n5678 & n5683;
  assign n5685 = n5684 ^ x32;
  assign n5745 = n5744 ^ n5685;
  assign n5675 = n5516 ^ n5450;
  assign n5676 = n5517 & n5675;
  assign n5677 = n5676 ^ n5450;
  assign n5746 = n5745 ^ n5677;
  assign n5667 = n1560 & n2527;
  assign n5668 = x81 & n2690;
  assign n5669 = x82 & n2530;
  assign n5670 = ~n5668 & ~n5669;
  assign n5671 = x83 & n2693;
  assign n5672 = n5670 & ~n5671;
  assign n5673 = ~n5667 & n5672;
  assign n5674 = n5673 ^ x29;
  assign n5747 = n5746 ^ n5674;
  assign n5664 = n5518 ^ n5439;
  assign n5665 = ~n5519 & ~n5664;
  assign n5666 = n5665 ^ n5439;
  assign n5748 = n5747 ^ n5666;
  assign n5656 = n1920 & n2102;
  assign n5657 = x84 & n2112;
  assign n5658 = x85 & n2105;
  assign n5659 = ~n5657 & ~n5658;
  assign n5660 = x86 & n2381;
  assign n5661 = n5659 & ~n5660;
  assign n5662 = ~n5656 & n5661;
  assign n5663 = n5662 ^ x26;
  assign n5749 = n5748 ^ n5663;
  assign n5653 = n5520 ^ n5428;
  assign n5654 = n5521 & n5653;
  assign n5655 = n5654 ^ n5428;
  assign n5750 = n5749 ^ n5655;
  assign n5645 = n1746 & n2310;
  assign n5646 = x88 & n1750;
  assign n5647 = x87 & n1871;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = x89 & n1873;
  assign n5650 = n5648 & ~n5649;
  assign n5651 = ~n5645 & n5650;
  assign n5652 = n5651 ^ x23;
  assign n5751 = n5750 ^ n5652;
  assign n5642 = n5522 ^ n5417;
  assign n5643 = ~n5523 & ~n5642;
  assign n5644 = n5643 ^ n5417;
  assign n5752 = n5751 ^ n5644;
  assign n5634 = n1404 & n2755;
  assign n5635 = x91 & n1408;
  assign n5636 = x90 & n1514;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = x92 & n1517;
  assign n5639 = n5637 & ~n5638;
  assign n5640 = ~n5634 & n5639;
  assign n5641 = n5640 ^ x20;
  assign n5753 = n5752 ^ n5641;
  assign n5631 = n5524 ^ n5406;
  assign n5632 = n5525 & n5631;
  assign n5633 = n5632 ^ n5406;
  assign n5754 = n5753 ^ n5633;
  assign n5623 = n1098 & n3247;
  assign n5624 = x94 & n1102;
  assign n5625 = x93 & n1198;
  assign n5626 = ~n5624 & ~n5625;
  assign n5627 = x95 & n1201;
  assign n5628 = n5626 & ~n5627;
  assign n5629 = ~n5623 & n5628;
  assign n5630 = n5629 ^ x17;
  assign n5755 = n5754 ^ n5630;
  assign n5620 = n5526 ^ n5395;
  assign n5621 = ~n5527 & ~n5620;
  assign n5622 = n5621 ^ n5395;
  assign n5756 = n5755 ^ n5622;
  assign n5612 = n821 & n3763;
  assign n5613 = x96 & n898;
  assign n5614 = x97 & n824;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = x98 & n901;
  assign n5617 = n5615 & ~n5616;
  assign n5618 = ~n5612 & n5617;
  assign n5619 = n5618 ^ x14;
  assign n5757 = n5756 ^ n5619;
  assign n5609 = n5528 ^ n5384;
  assign n5610 = n5529 & n5609;
  assign n5611 = n5610 ^ n5384;
  assign n5758 = n5757 ^ n5611;
  assign n5601 = n596 & n4323;
  assign n5602 = x99 & n673;
  assign n5603 = x101 & n676;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = x100 & n601;
  assign n5606 = n5604 & ~n5605;
  assign n5607 = ~n5601 & n5606;
  assign n5608 = n5607 ^ x11;
  assign n5759 = n5758 ^ n5608;
  assign n5598 = n5530 ^ n5373;
  assign n5599 = ~n5531 & ~n5598;
  assign n5600 = n5599 ^ n5373;
  assign n5760 = n5759 ^ n5600;
  assign n5590 = n399 & n4912;
  assign n5591 = x102 & n478;
  assign n5592 = x103 & n402;
  assign n5593 = ~n5591 & ~n5592;
  assign n5594 = x104 & n470;
  assign n5595 = n5593 & ~n5594;
  assign n5596 = ~n5590 & n5595;
  assign n5597 = n5596 ^ x8;
  assign n5761 = n5760 ^ n5597;
  assign n5587 = n5532 ^ n5362;
  assign n5588 = n5533 & n5587;
  assign n5589 = n5588 ^ n5362;
  assign n5762 = n5761 ^ n5589;
  assign n5578 = n4896 ^ x107;
  assign n5579 = n239 & n5578;
  assign n5580 = x105 & n249;
  assign n5581 = x107 & n280;
  assign n5582 = ~n5580 & ~n5581;
  assign n5583 = x106 & n242;
  assign n5584 = n5582 & ~n5583;
  assign n5585 = ~n5579 & n5584;
  assign n5586 = n5585 ^ x5;
  assign n5763 = n5762 ^ n5586;
  assign n5575 = n5534 ^ n5350;
  assign n5576 = ~n5535 & n5575;
  assign n5577 = n5576 ^ n5350;
  assign n5764 = n5763 ^ n5577;
  assign n5554 = x109 ^ x108;
  assign n5555 = n5554 ^ n5335;
  assign n5556 = n4894 ^ x109;
  assign n5557 = n5556 ^ n4894;
  assign n5558 = n5336 & ~n5557;
  assign n5559 = n5558 ^ n4894;
  assign n5560 = n5559 ^ n5554;
  assign n5561 = n5555 & ~n5560;
  assign n5562 = n5561 ^ n5558;
  assign n5563 = n5562 ^ n4894;
  assign n5564 = n5563 ^ n5335;
  assign n5565 = n5554 & ~n5564;
  assign n5566 = n5565 ^ n5554;
  assign n5567 = n5566 ^ x108;
  assign n5568 = n5567 ^ x109;
  assign n5569 = n169 & ~n5568;
  assign n5570 = n5569 ^ x1;
  assign n5571 = n5570 ^ x110;
  assign n5542 = x109 ^ x2;
  assign n5543 = n5542 ^ x1;
  assign n5544 = n5543 ^ n5542;
  assign n5545 = n5544 ^ x0;
  assign n5546 = n5542 ^ x109;
  assign n5547 = n5546 ^ x108;
  assign n5548 = ~x108 & ~n5547;
  assign n5549 = n5548 ^ n5542;
  assign n5550 = n5549 ^ x108;
  assign n5551 = n5545 & ~n5550;
  assign n5552 = n5551 ^ n5548;
  assign n5553 = n5552 ^ x108;
  assign n5572 = n5571 ^ n5553;
  assign n5573 = ~x0 & ~n5572;
  assign n5574 = n5573 ^ n5571;
  assign n5765 = n5764 ^ n5574;
  assign n5539 = n5536 ^ n5322;
  assign n5540 = n5537 & ~n5539;
  assign n5541 = n5540 ^ n5322;
  assign n5766 = n5765 ^ n5541;
  assign n5970 = n5715 ^ n5704;
  assign n5971 = n5713 & ~n5970;
  assign n5972 = n5971 ^ n5715;
  assign n5941 = x47 ^ x46;
  assign n5942 = n5481 & n5941;
  assign n5943 = n142 & n5942;
  assign n5944 = ~x44 & ~x45;
  assign n5945 = n5944 ^ n5709;
  assign n5946 = x46 & n5945;
  assign n5947 = n5946 ^ n5709;
  assign n5948 = ~n5943 & ~n5947;
  assign n5949 = x65 & ~n5948;
  assign n5950 = n152 & n5941;
  assign n5951 = x66 & n5481;
  assign n5952 = ~n5950 & n5951;
  assign n5953 = ~n5949 & ~n5952;
  assign n5962 = ~x46 & x47;
  assign n5963 = n5944 & n5962;
  assign n5964 = x64 & n5963;
  assign n5965 = n5953 & ~n5964;
  assign n5957 = x46 ^ x44;
  assign n5958 = x64 & n5957;
  assign n5959 = n5958 ^ n233;
  assign n5960 = ~n5481 & ~n5959;
  assign n5961 = n5960 ^ n233;
  assign n5966 = n5965 ^ n5961;
  assign n5954 = x46 & x64;
  assign n5955 = n5709 & n5954;
  assign n5956 = n5953 & ~n5955;
  assign n5967 = n5966 ^ n5956;
  assign n5968 = ~x47 & ~n5967;
  assign n5969 = n5968 ^ n5966;
  assign n5973 = n5972 ^ n5969;
  assign n5933 = n420 & n5262;
  assign n5934 = x68 & n5266;
  assign n5935 = x67 & n5488;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = x69 & n5491;
  assign n5938 = n5936 & ~n5937;
  assign n5939 = ~n5933 & n5938;
  assign n5940 = n5939 ^ x44;
  assign n5974 = n5973 ^ n5940;
  assign n5930 = n5727 ^ n5716;
  assign n5931 = ~n5728 & ~n5930;
  assign n5932 = n5931 ^ n5719;
  assign n5975 = n5974 ^ n5932;
  assign n5922 = n575 & n4643;
  assign n5923 = x71 & n4646;
  assign n5924 = x70 & n4653;
  assign n5925 = ~n5923 & ~n5924;
  assign n5926 = x72 & n5046;
  assign n5927 = n5925 & ~n5926;
  assign n5928 = ~n5922 & n5927;
  assign n5929 = n5928 ^ x41;
  assign n5976 = n5975 ^ n5929;
  assign n5919 = n5729 ^ n5688;
  assign n5920 = n5730 & n5919;
  assign n5921 = n5920 ^ n5688;
  assign n5977 = n5976 ^ n5921;
  assign n5911 = n789 & n4040;
  assign n5912 = x74 & n4044;
  assign n5913 = x75 & n4270;
  assign n5914 = ~n5912 & ~n5913;
  assign n5915 = x73 & n4267;
  assign n5916 = n5914 & ~n5915;
  assign n5917 = ~n5911 & n5916;
  assign n5918 = n5917 ^ x38;
  assign n5978 = n5977 ^ n5918;
  assign n5903 = n1041 & n3522;
  assign n5904 = x76 & n3699;
  assign n5905 = x78 & n3701;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = x77 & n3526;
  assign n5908 = n5906 & ~n5907;
  assign n5909 = ~n5903 & n5908;
  assign n5910 = n5909 ^ x35;
  assign n5979 = n5978 ^ n5910;
  assign n5900 = n5742 ^ n5731;
  assign n5901 = ~n5743 & ~n5900;
  assign n5902 = n5901 ^ n5734;
  assign n5980 = n5979 ^ n5902;
  assign n5892 = n1340 & n3009;
  assign n5893 = x79 & n3181;
  assign n5894 = x80 & n3013;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = x81 & n3183;
  assign n5897 = n5895 & ~n5896;
  assign n5898 = ~n5892 & n5897;
  assign n5899 = n5898 ^ x32;
  assign n5981 = n5980 ^ n5899;
  assign n5889 = n5744 ^ n5677;
  assign n5890 = n5745 & n5889;
  assign n5891 = n5890 ^ n5677;
  assign n5982 = n5981 ^ n5891;
  assign n5881 = n1667 & n2527;
  assign n5882 = x83 & n2530;
  assign n5883 = x82 & n2690;
  assign n5884 = ~n5882 & ~n5883;
  assign n5885 = x84 & n2693;
  assign n5886 = n5884 & ~n5885;
  assign n5887 = ~n5881 & n5886;
  assign n5888 = n5887 ^ x29;
  assign n5983 = n5982 ^ n5888;
  assign n5878 = n5746 ^ n5666;
  assign n5879 = ~n5747 & ~n5878;
  assign n5880 = n5879 ^ n5666;
  assign n5984 = n5983 ^ n5880;
  assign n5870 = n2039 & n2102;
  assign n5871 = x85 & n2112;
  assign n5872 = x86 & n2105;
  assign n5873 = ~n5871 & ~n5872;
  assign n5874 = x87 & n2381;
  assign n5875 = n5873 & ~n5874;
  assign n5876 = ~n5870 & n5875;
  assign n5877 = n5876 ^ x26;
  assign n5985 = n5984 ^ n5877;
  assign n5867 = n5748 ^ n5655;
  assign n5868 = n5749 & n5867;
  assign n5869 = n5868 ^ n5655;
  assign n5986 = n5985 ^ n5869;
  assign n5859 = n1746 & n2448;
  assign n5860 = x89 & n1750;
  assign n5861 = x88 & n1871;
  assign n5862 = ~n5860 & ~n5861;
  assign n5863 = x90 & n1873;
  assign n5864 = n5862 & ~n5863;
  assign n5865 = ~n5859 & n5864;
  assign n5866 = n5865 ^ x23;
  assign n5987 = n5986 ^ n5866;
  assign n5856 = n5750 ^ n5644;
  assign n5857 = ~n5751 & ~n5856;
  assign n5858 = n5857 ^ n5644;
  assign n5988 = n5987 ^ n5858;
  assign n5848 = n1404 & n2901;
  assign n5849 = x92 & n1408;
  assign n5850 = x91 & n1514;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = x93 & n1517;
  assign n5853 = n5851 & ~n5852;
  assign n5854 = ~n5848 & n5853;
  assign n5855 = n5854 ^ x20;
  assign n5989 = n5988 ^ n5855;
  assign n5845 = n5752 ^ n5633;
  assign n5846 = n5753 & n5845;
  assign n5847 = n5846 ^ n5633;
  assign n5990 = n5989 ^ n5847;
  assign n5837 = n1098 & n3403;
  assign n5838 = x94 & n1198;
  assign n5839 = x95 & n1102;
  assign n5840 = ~n5838 & ~n5839;
  assign n5841 = x96 & n1201;
  assign n5842 = n5840 & ~n5841;
  assign n5843 = ~n5837 & n5842;
  assign n5844 = n5843 ^ x17;
  assign n5991 = n5990 ^ n5844;
  assign n5834 = n5754 ^ n5622;
  assign n5835 = ~n5755 & ~n5834;
  assign n5836 = n5835 ^ n5622;
  assign n5992 = n5991 ^ n5836;
  assign n5826 = n821 & n3943;
  assign n5827 = x97 & n898;
  assign n5828 = x98 & n824;
  assign n5829 = ~n5827 & ~n5828;
  assign n5830 = x99 & n901;
  assign n5831 = n5829 & ~n5830;
  assign n5832 = ~n5826 & n5831;
  assign n5833 = n5832 ^ x14;
  assign n5993 = n5992 ^ n5833;
  assign n5823 = n5756 ^ n5611;
  assign n5824 = n5757 & n5823;
  assign n5825 = n5824 ^ n5611;
  assign n5994 = n5993 ^ n5825;
  assign n5815 = n596 & n4509;
  assign n5816 = x100 & n673;
  assign n5817 = x101 & n601;
  assign n5818 = ~n5816 & ~n5817;
  assign n5819 = x102 & n676;
  assign n5820 = n5818 & ~n5819;
  assign n5821 = ~n5815 & n5820;
  assign n5822 = n5821 ^ x11;
  assign n5995 = n5994 ^ n5822;
  assign n5812 = n5758 ^ n5600;
  assign n5813 = ~n5759 & ~n5812;
  assign n5814 = n5813 ^ n5600;
  assign n5996 = n5995 ^ n5814;
  assign n5804 = n399 & n5117;
  assign n5805 = x103 & n478;
  assign n5806 = x104 & n402;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = x105 & n470;
  assign n5809 = n5807 & ~n5808;
  assign n5810 = ~n5804 & n5809;
  assign n5811 = n5810 ^ x8;
  assign n5997 = n5996 ^ n5811;
  assign n5801 = n5760 ^ n5589;
  assign n5802 = n5761 & n5801;
  assign n5803 = n5802 ^ n5589;
  assign n5998 = n5997 ^ n5803;
  assign n5792 = n5107 ^ x108;
  assign n5793 = n239 & n5792;
  assign n5794 = x106 & n249;
  assign n5795 = x108 & n280;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = x107 & n242;
  assign n5798 = n5796 & ~n5797;
  assign n5799 = ~n5793 & n5798;
  assign n5800 = n5799 ^ x5;
  assign n5999 = n5998 ^ n5800;
  assign n5789 = n5762 ^ n5577;
  assign n5790 = ~n5763 & n5789;
  assign n5791 = n5790 ^ n5577;
  assign n6000 = n5999 ^ n5791;
  assign n5778 = x109 & n5567;
  assign n5779 = ~x110 & ~n5778;
  assign n5780 = ~x109 & ~n5567;
  assign n5781 = x110 & ~n5780;
  assign n5782 = ~n5779 & ~n5781;
  assign n5783 = n169 & ~n5782;
  assign n5784 = n5783 ^ x1;
  assign n5785 = n5784 ^ x111;
  assign n5770 = x110 ^ x2;
  assign n5771 = n5770 ^ x109;
  assign n5772 = n5771 ^ n5770;
  assign n5773 = n5770 ^ x110;
  assign n5774 = ~n5772 & n5773;
  assign n5775 = n5774 ^ n5770;
  assign n5776 = ~x1 & n5775;
  assign n5777 = n5776 ^ n5770;
  assign n5786 = n5785 ^ n5777;
  assign n5787 = ~x0 & n5786;
  assign n5788 = n5787 ^ n5785;
  assign n6001 = n6000 ^ n5788;
  assign n5767 = n5764 ^ n5541;
  assign n5768 = n5765 & ~n5767;
  assign n5769 = n5768 ^ n5541;
  assign n6002 = n6001 ^ n5769;
  assign n6193 = n5961 & n5965;
  assign n6194 = x47 & n6193;
  assign n6191 = x48 ^ x47;
  assign n6192 = x64 & n6191;
  assign n6195 = n6194 ^ n6192;
  assign n6178 = n168 & n5941;
  assign n6179 = n6178 ^ x67;
  assign n6180 = n5481 & n6179;
  assign n6181 = x66 & n5947;
  assign n6182 = n5709 ^ x47;
  assign n6183 = n6182 ^ n5709;
  assign n6184 = n5945 & n6183;
  assign n6185 = n6184 ^ n5709;
  assign n6186 = n5941 & n6185;
  assign n6187 = x65 & n6186;
  assign n6188 = ~n6181 & ~n6187;
  assign n6189 = ~n6180 & n6188;
  assign n6190 = n6189 ^ x47;
  assign n6196 = n6195 ^ n6190;
  assign n6170 = n458 & n5262;
  assign n6171 = x69 & n5266;
  assign n6172 = x68 & n5488;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = x70 & n5491;
  assign n6175 = n6173 & ~n6174;
  assign n6176 = ~n6170 & n6175;
  assign n6177 = n6176 ^ x44;
  assign n6197 = n6196 ^ n6177;
  assign n6167 = n5969 ^ n5940;
  assign n6168 = n5973 & n6167;
  assign n6169 = n6168 ^ n5972;
  assign n6198 = n6197 ^ n6169;
  assign n6164 = n5974 ^ n5929;
  assign n6165 = ~n5975 & ~n6164;
  assign n6166 = n6165 ^ n5932;
  assign n6199 = n6198 ^ n6166;
  assign n6156 = ~n653 & n4643;
  assign n6157 = x72 & n4646;
  assign n6158 = x71 & n4653;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = x73 & n5046;
  assign n6161 = n6159 & ~n6160;
  assign n6162 = ~n6156 & n6161;
  assign n6163 = n6162 ^ x41;
  assign n6200 = n6199 ^ n6163;
  assign n6148 = n870 & n4040;
  assign n6149 = x74 & n4267;
  assign n6150 = x76 & n4270;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = x75 & n4044;
  assign n6153 = n6151 & ~n6152;
  assign n6154 = ~n6148 & n6153;
  assign n6155 = n6154 ^ x38;
  assign n6201 = n6200 ^ n6155;
  assign n6145 = n5976 ^ n5918;
  assign n6146 = n5977 & n6145;
  assign n6147 = n6146 ^ n5921;
  assign n6202 = n6201 ^ n6147;
  assign n6142 = n5978 ^ n5902;
  assign n6143 = ~n5979 & ~n6142;
  assign n6144 = n6143 ^ n5902;
  assign n6203 = n6202 ^ n6144;
  assign n6134 = n1149 & n3522;
  assign n6135 = x77 & n3699;
  assign n6136 = x78 & n3526;
  assign n6137 = ~n6135 & ~n6136;
  assign n6138 = x79 & n3701;
  assign n6139 = n6137 & ~n6138;
  assign n6140 = ~n6134 & n6139;
  assign n6141 = n6140 ^ x35;
  assign n6204 = n6203 ^ n6141;
  assign n6126 = n1454 & n3009;
  assign n6127 = x80 & n3181;
  assign n6128 = x81 & n3013;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = x82 & n3183;
  assign n6131 = n6129 & ~n6130;
  assign n6132 = ~n6126 & n6131;
  assign n6133 = n6132 ^ x32;
  assign n6205 = n6204 ^ n6133;
  assign n6123 = n5980 ^ n5891;
  assign n6124 = n5981 & n6123;
  assign n6125 = n6124 ^ n5891;
  assign n6206 = n6205 ^ n6125;
  assign n6115 = n1801 & n2527;
  assign n6116 = x84 & n2530;
  assign n6117 = x83 & n2690;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = x85 & n2693;
  assign n6120 = n6118 & ~n6119;
  assign n6121 = ~n6115 & n6120;
  assign n6122 = n6121 ^ x29;
  assign n6207 = n6206 ^ n6122;
  assign n6112 = n5982 ^ n5880;
  assign n6113 = ~n5983 & ~n6112;
  assign n6114 = n6113 ^ n5880;
  assign n6208 = n6207 ^ n6114;
  assign n6104 = n2102 & n2176;
  assign n6105 = x87 & n2105;
  assign n6106 = x86 & n2112;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = x88 & n2381;
  assign n6109 = n6107 & ~n6108;
  assign n6110 = ~n6104 & n6109;
  assign n6111 = n6110 ^ x26;
  assign n6209 = n6208 ^ n6111;
  assign n6101 = n5984 ^ n5869;
  assign n6102 = n5985 & n6101;
  assign n6103 = n6102 ^ n5869;
  assign n6210 = n6209 ^ n6103;
  assign n6093 = n1746 & n2607;
  assign n6094 = x89 & n1871;
  assign n6095 = x90 & n1750;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = x91 & n1873;
  assign n6098 = n6096 & ~n6097;
  assign n6099 = ~n6093 & n6098;
  assign n6100 = n6099 ^ x23;
  assign n6211 = n6210 ^ n6100;
  assign n6090 = n5986 ^ n5858;
  assign n6091 = ~n5987 & ~n6090;
  assign n6092 = n6091 ^ n5858;
  assign n6212 = n6211 ^ n6092;
  assign n6082 = n1404 & n3078;
  assign n6083 = x93 & n1408;
  assign n6084 = x92 & n1514;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = x94 & n1517;
  assign n6087 = n6085 & ~n6086;
  assign n6088 = ~n6082 & n6087;
  assign n6089 = n6088 ^ x20;
  assign n6213 = n6212 ^ n6089;
  assign n6079 = n5988 ^ n5847;
  assign n6080 = n5989 & n6079;
  assign n6081 = n6080 ^ n5847;
  assign n6214 = n6213 ^ n6081;
  assign n6071 = n1098 & n3585;
  assign n6072 = x96 & n1102;
  assign n6073 = x95 & n1198;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = x97 & n1201;
  assign n6076 = n6074 & ~n6075;
  assign n6077 = ~n6071 & n6076;
  assign n6078 = n6077 ^ x17;
  assign n6215 = n6214 ^ n6078;
  assign n6068 = n5990 ^ n5836;
  assign n6069 = ~n5991 & ~n6068;
  assign n6070 = n6069 ^ n5836;
  assign n6216 = n6215 ^ n6070;
  assign n6060 = n821 & n4141;
  assign n6061 = x98 & n898;
  assign n6062 = x100 & n901;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = x99 & n824;
  assign n6065 = n6063 & ~n6064;
  assign n6066 = ~n6060 & n6065;
  assign n6067 = n6066 ^ x14;
  assign n6217 = n6216 ^ n6067;
  assign n6057 = n5992 ^ n5825;
  assign n6058 = n5993 & n6057;
  assign n6059 = n6058 ^ n5825;
  assign n6218 = n6217 ^ n6059;
  assign n6049 = n596 & n4718;
  assign n6050 = x101 & n673;
  assign n6051 = x103 & n676;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = x102 & n601;
  assign n6054 = n6052 & ~n6053;
  assign n6055 = ~n6049 & n6054;
  assign n6056 = n6055 ^ x11;
  assign n6219 = n6218 ^ n6056;
  assign n6046 = n5994 ^ n5814;
  assign n6047 = ~n5995 & ~n6046;
  assign n6048 = n6047 ^ n5814;
  assign n6220 = n6219 ^ n6048;
  assign n6038 = n399 & n5351;
  assign n6039 = x104 & n478;
  assign n6040 = x105 & n402;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = x106 & n470;
  assign n6043 = n6041 & ~n6042;
  assign n6044 = ~n6038 & n6043;
  assign n6045 = n6044 ^ x8;
  assign n6221 = n6220 ^ n6045;
  assign n6035 = n5996 ^ n5803;
  assign n6036 = n5997 & n6035;
  assign n6037 = n6036 ^ n5803;
  assign n6222 = n6221 ^ n6037;
  assign n6026 = n5341 ^ x109;
  assign n6027 = n239 & n6026;
  assign n6028 = x107 & n249;
  assign n6029 = x108 & n242;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = x109 & n280;
  assign n6032 = n6030 & ~n6031;
  assign n6033 = ~n6027 & n6032;
  assign n6034 = n6033 ^ x5;
  assign n6223 = n6222 ^ n6034;
  assign n6023 = n5998 ^ n5791;
  assign n6024 = ~n5999 & n6023;
  assign n6025 = n6024 ^ n5791;
  assign n6224 = n6223 ^ n6025;
  assign n6012 = x111 ^ x2;
  assign n6013 = n6012 ^ x110;
  assign n6014 = n6013 ^ n6012;
  assign n6015 = n6012 ^ x111;
  assign n6016 = ~n6014 & n6015;
  assign n6017 = n6016 ^ n6012;
  assign n6018 = ~x1 & n6017;
  assign n6019 = n6018 ^ n6012;
  assign n6006 = ~x111 & ~n5781;
  assign n6007 = x111 & ~n5779;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = n169 & ~n6008;
  assign n6010 = n6009 ^ x1;
  assign n6011 = n6010 ^ x112;
  assign n6020 = n6019 ^ n6011;
  assign n6021 = ~x0 & n6020;
  assign n6022 = n6021 ^ n6011;
  assign n6225 = n6224 ^ n6022;
  assign n6003 = n6000 ^ n5769;
  assign n6004 = n6001 & ~n6003;
  assign n6005 = n6004 ^ n5769;
  assign n6226 = n6225 ^ n6005;
  assign n6419 = ~n6192 & ~n6194;
  assign n6420 = ~n6190 & ~n6419;
  assign n6414 = x65 ^ x48;
  assign n6415 = n6191 & ~n6414;
  assign n6416 = n6415 ^ x47;
  assign n6417 = n6416 ^ x49;
  assign n6411 = x47 & x48;
  assign n6412 = n6411 ^ x49;
  assign n6413 = ~x64 & n6412;
  assign n6418 = n6417 ^ n6413;
  assign n6421 = n6420 ^ n6418;
  assign n6402 = n321 & n5942;
  assign n6403 = x66 & n6186;
  assign n6404 = x67 & n5947;
  assign n6405 = ~n6403 & ~n6404;
  assign n6406 = n5481 & ~n5941;
  assign n6407 = x68 & n6406;
  assign n6408 = n6405 & ~n6407;
  assign n6409 = ~n6402 & n6408;
  assign n6410 = n6409 ^ x47;
  assign n6422 = n6421 ^ n6410;
  assign n6394 = n517 & n5262;
  assign n6395 = x69 & n5488;
  assign n6396 = x70 & n5266;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = x71 & n5491;
  assign n6399 = n6397 & ~n6398;
  assign n6400 = ~n6394 & n6399;
  assign n6401 = n6400 ^ x44;
  assign n6423 = n6422 ^ n6401;
  assign n6391 = n6196 ^ n6169;
  assign n6392 = ~n6197 & ~n6391;
  assign n6393 = n6392 ^ n6169;
  assign n6424 = n6423 ^ n6393;
  assign n6383 = ~n721 & n4643;
  assign n6384 = x73 & n4646;
  assign n6385 = x72 & n4653;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = x74 & n5046;
  assign n6388 = n6386 & ~n6387;
  assign n6389 = ~n6383 & n6388;
  assign n6390 = n6389 ^ x41;
  assign n6425 = n6424 ^ n6390;
  assign n6380 = n6198 ^ n6163;
  assign n6381 = n6199 & n6380;
  assign n6382 = n6381 ^ n6166;
  assign n6426 = n6425 ^ n6382;
  assign n6372 = n956 & n4040;
  assign n6373 = x75 & n4267;
  assign n6374 = x76 & n4044;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = x77 & n4270;
  assign n6377 = n6375 & ~n6376;
  assign n6378 = ~n6372 & n6377;
  assign n6379 = n6378 ^ x38;
  assign n6427 = n6426 ^ n6379;
  assign n6369 = n6200 ^ n6147;
  assign n6370 = ~n6201 & ~n6369;
  assign n6371 = n6370 ^ n6147;
  assign n6428 = n6427 ^ n6371;
  assign n6361 = n1242 & n3522;
  assign n6362 = x78 & n3699;
  assign n6363 = x79 & n3526;
  assign n6364 = ~n6362 & ~n6363;
  assign n6365 = x80 & n3701;
  assign n6366 = n6364 & ~n6365;
  assign n6367 = ~n6361 & n6366;
  assign n6368 = n6367 ^ x35;
  assign n6429 = n6428 ^ n6368;
  assign n6358 = n6202 ^ n6141;
  assign n6359 = n6203 & n6358;
  assign n6360 = n6359 ^ n6144;
  assign n6430 = n6429 ^ n6360;
  assign n6350 = n1560 & n3009;
  assign n6351 = x81 & n3181;
  assign n6352 = x82 & n3013;
  assign n6353 = ~n6351 & ~n6352;
  assign n6354 = x83 & n3183;
  assign n6355 = n6353 & ~n6354;
  assign n6356 = ~n6350 & n6355;
  assign n6357 = n6356 ^ x32;
  assign n6431 = n6430 ^ n6357;
  assign n6347 = n6204 ^ n6125;
  assign n6348 = ~n6205 & ~n6347;
  assign n6349 = n6348 ^ n6125;
  assign n6432 = n6431 ^ n6349;
  assign n6339 = n1920 & n2527;
  assign n6340 = x84 & n2690;
  assign n6341 = x85 & n2530;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = x86 & n2693;
  assign n6344 = n6342 & ~n6343;
  assign n6345 = ~n6339 & n6344;
  assign n6346 = n6345 ^ x29;
  assign n6433 = n6432 ^ n6346;
  assign n6336 = n6206 ^ n6114;
  assign n6337 = n6207 & n6336;
  assign n6338 = n6337 ^ n6114;
  assign n6434 = n6433 ^ n6338;
  assign n6328 = n2102 & n2310;
  assign n6329 = x87 & n2112;
  assign n6330 = x88 & n2105;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = x89 & n2381;
  assign n6333 = n6331 & ~n6332;
  assign n6334 = ~n6328 & n6333;
  assign n6335 = n6334 ^ x26;
  assign n6435 = n6434 ^ n6335;
  assign n6325 = n6208 ^ n6103;
  assign n6326 = ~n6209 & ~n6325;
  assign n6327 = n6326 ^ n6103;
  assign n6436 = n6435 ^ n6327;
  assign n6317 = n1746 & n2755;
  assign n6318 = x91 & n1750;
  assign n6319 = x90 & n1871;
  assign n6320 = ~n6318 & ~n6319;
  assign n6321 = x92 & n1873;
  assign n6322 = n6320 & ~n6321;
  assign n6323 = ~n6317 & n6322;
  assign n6324 = n6323 ^ x23;
  assign n6437 = n6436 ^ n6324;
  assign n6314 = n6210 ^ n6092;
  assign n6315 = n6211 & n6314;
  assign n6316 = n6315 ^ n6092;
  assign n6438 = n6437 ^ n6316;
  assign n6306 = n1404 & n3247;
  assign n6307 = x93 & n1514;
  assign n6308 = x94 & n1408;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = x95 & n1517;
  assign n6311 = n6309 & ~n6310;
  assign n6312 = ~n6306 & n6311;
  assign n6313 = n6312 ^ x20;
  assign n6439 = n6438 ^ n6313;
  assign n6303 = n6212 ^ n6081;
  assign n6304 = ~n6213 & ~n6303;
  assign n6305 = n6304 ^ n6081;
  assign n6440 = n6439 ^ n6305;
  assign n6295 = n1098 & n3763;
  assign n6296 = x97 & n1102;
  assign n6297 = x96 & n1198;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = x98 & n1201;
  assign n6300 = n6298 & ~n6299;
  assign n6301 = ~n6295 & n6300;
  assign n6302 = n6301 ^ x17;
  assign n6441 = n6440 ^ n6302;
  assign n6292 = n6214 ^ n6070;
  assign n6293 = n6215 & n6292;
  assign n6294 = n6293 ^ n6070;
  assign n6442 = n6441 ^ n6294;
  assign n6284 = n821 & n4323;
  assign n6285 = x99 & n898;
  assign n6286 = x100 & n824;
  assign n6287 = ~n6285 & ~n6286;
  assign n6288 = x101 & n901;
  assign n6289 = n6287 & ~n6288;
  assign n6290 = ~n6284 & n6289;
  assign n6291 = n6290 ^ x14;
  assign n6443 = n6442 ^ n6291;
  assign n6281 = n6216 ^ n6059;
  assign n6282 = ~n6217 & ~n6281;
  assign n6283 = n6282 ^ n6059;
  assign n6444 = n6443 ^ n6283;
  assign n6273 = n596 & n4912;
  assign n6274 = x102 & n673;
  assign n6275 = x103 & n601;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = x104 & n676;
  assign n6278 = n6276 & ~n6277;
  assign n6279 = ~n6273 & n6278;
  assign n6280 = n6279 ^ x11;
  assign n6445 = n6444 ^ n6280;
  assign n6270 = n6218 ^ n6048;
  assign n6271 = n6219 & n6270;
  assign n6272 = n6271 ^ n6048;
  assign n6446 = n6445 ^ n6272;
  assign n6262 = n399 & n5578;
  assign n6263 = x105 & n478;
  assign n6264 = x106 & n402;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = x107 & n470;
  assign n6267 = n6265 & ~n6266;
  assign n6268 = ~n6262 & n6267;
  assign n6269 = n6268 ^ x8;
  assign n6447 = n6446 ^ n6269;
  assign n6259 = n6220 ^ n6037;
  assign n6260 = ~n6221 & ~n6259;
  assign n6261 = n6260 ^ n6037;
  assign n6448 = n6447 ^ n6261;
  assign n6249 = x110 ^ x109;
  assign n6250 = n6249 ^ n5567;
  assign n6251 = n239 & n6250;
  assign n6252 = x108 & n249;
  assign n6253 = x109 & n242;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = x110 & n280;
  assign n6256 = n6254 & ~n6255;
  assign n6257 = ~n6251 & n6256;
  assign n6258 = n6257 ^ x5;
  assign n6449 = n6448 ^ n6258;
  assign n6246 = n6222 ^ n6025;
  assign n6247 = n6223 & ~n6246;
  assign n6248 = n6247 ^ n6025;
  assign n6450 = n6449 ^ n6248;
  assign n6232 = x112 ^ x111;
  assign n6233 = ~n6008 & n6232;
  assign n6234 = n169 & ~n6233;
  assign n6235 = n6234 ^ x1;
  assign n6236 = n6235 ^ x113;
  assign n6230 = x1 & x112;
  assign n6231 = n6230 ^ x2;
  assign n6237 = n6236 ^ n6231;
  assign n6238 = n6237 ^ n6236;
  assign n6239 = x111 & n197;
  assign n6240 = n6239 ^ n6236;
  assign n6241 = n6240 ^ n6236;
  assign n6242 = n6238 & ~n6241;
  assign n6243 = n6242 ^ n6236;
  assign n6244 = ~x0 & n6243;
  assign n6245 = n6244 ^ n6236;
  assign n6451 = n6450 ^ n6245;
  assign n6227 = n6224 ^ n6005;
  assign n6228 = ~n6225 & n6227;
  assign n6229 = n6228 ^ n6005;
  assign n6452 = n6451 ^ n6229;
  assign n6670 = n789 & n4643;
  assign n6671 = x73 & n4653;
  assign n6672 = x75 & n5046;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = x74 & n4646;
  assign n6675 = n6673 & ~n6674;
  assign n6676 = ~n6670 & n6675;
  assign n6677 = n6676 ^ x41;
  assign n6667 = n6424 ^ n6382;
  assign n6668 = n6425 & n6667;
  assign n6669 = n6668 ^ n6382;
  assign n6678 = n6677 ^ n6669;
  assign n6654 = n420 & n5942;
  assign n6655 = x68 & n5947;
  assign n6656 = x67 & n6186;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = x69 & n6406;
  assign n6659 = n6657 & ~n6658;
  assign n6660 = ~n6654 & n6659;
  assign n6661 = n6660 ^ x47;
  assign n6622 = ~x47 & ~x48;
  assign n6644 = ~n233 & ~n6622;
  assign n6645 = n6644 ^ n6411;
  assign n6646 = x64 ^ x49;
  assign n6647 = n6646 ^ x49;
  assign n6648 = n6644 ^ x49;
  assign n6649 = ~n6647 & n6648;
  assign n6650 = n6649 ^ x49;
  assign n6651 = ~n6645 & ~n6650;
  assign n6652 = n6651 ^ n6411;
  assign n6653 = x50 & n6652;
  assign n6662 = n6661 ^ n6653;
  assign n6623 = ~x49 & x64;
  assign n6624 = n6622 & n6623;
  assign n6625 = x50 ^ x49;
  assign n6626 = n6191 & n6625;
  assign n6627 = n142 & n6626;
  assign n6628 = n6622 ^ n6411;
  assign n6629 = x49 & n6628;
  assign n6630 = n6629 ^ n6411;
  assign n6631 = ~n6627 & ~n6630;
  assign n6632 = x65 & ~n6631;
  assign n6633 = n152 & n6625;
  assign n6634 = x66 & n6191;
  assign n6635 = ~n6633 & n6634;
  assign n6636 = ~n6632 & ~n6635;
  assign n6637 = n6636 ^ x50;
  assign n6638 = x49 & x64;
  assign n6639 = n6411 & n6638;
  assign n6640 = n6636 & n6639;
  assign n6641 = n6637 & n6640;
  assign n6642 = n6641 ^ n6637;
  assign n6643 = ~n6624 & ~n6642;
  assign n6663 = n6662 ^ n6643;
  assign n6619 = n6418 ^ n6410;
  assign n6620 = n6421 & n6619;
  assign n6621 = n6620 ^ n6420;
  assign n6664 = n6663 ^ n6621;
  assign n6616 = n6422 ^ n6393;
  assign n6617 = ~n6423 & ~n6616;
  assign n6618 = n6617 ^ n6393;
  assign n6665 = n6664 ^ n6618;
  assign n6608 = n575 & n5262;
  assign n6609 = x71 & n5266;
  assign n6610 = x70 & n5488;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = x72 & n5491;
  assign n6613 = n6611 & ~n6612;
  assign n6614 = ~n6608 & n6613;
  assign n6615 = n6614 ^ x44;
  assign n6666 = n6665 ^ n6615;
  assign n6679 = n6678 ^ n6666;
  assign n6600 = n1041 & n4040;
  assign n6601 = x76 & n4267;
  assign n6602 = x78 & n4270;
  assign n6603 = ~n6601 & ~n6602;
  assign n6604 = x77 & n4044;
  assign n6605 = n6603 & ~n6604;
  assign n6606 = ~n6600 & n6605;
  assign n6607 = n6606 ^ x38;
  assign n6680 = n6679 ^ n6607;
  assign n6597 = n6426 ^ n6371;
  assign n6598 = ~n6427 & ~n6597;
  assign n6599 = n6598 ^ n6371;
  assign n6681 = n6680 ^ n6599;
  assign n6589 = n1340 & n3522;
  assign n6590 = x79 & n3699;
  assign n6591 = x81 & n3701;
  assign n6592 = ~n6590 & ~n6591;
  assign n6593 = x80 & n3526;
  assign n6594 = n6592 & ~n6593;
  assign n6595 = ~n6589 & n6594;
  assign n6596 = n6595 ^ x35;
  assign n6682 = n6681 ^ n6596;
  assign n6586 = n6428 ^ n6360;
  assign n6587 = n6429 & n6586;
  assign n6588 = n6587 ^ n6360;
  assign n6683 = n6682 ^ n6588;
  assign n6578 = n1667 & n3009;
  assign n6579 = x83 & n3013;
  assign n6580 = x82 & n3181;
  assign n6581 = ~n6579 & ~n6580;
  assign n6582 = x84 & n3183;
  assign n6583 = n6581 & ~n6582;
  assign n6584 = ~n6578 & n6583;
  assign n6585 = n6584 ^ x32;
  assign n6684 = n6683 ^ n6585;
  assign n6575 = n6430 ^ n6349;
  assign n6576 = ~n6431 & ~n6575;
  assign n6577 = n6576 ^ n6349;
  assign n6685 = n6684 ^ n6577;
  assign n6567 = n2039 & n2527;
  assign n6568 = x85 & n2690;
  assign n6569 = x86 & n2530;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = x87 & n2693;
  assign n6572 = n6570 & ~n6571;
  assign n6573 = ~n6567 & n6572;
  assign n6574 = n6573 ^ x29;
  assign n6686 = n6685 ^ n6574;
  assign n6564 = n6432 ^ n6338;
  assign n6565 = n6433 & n6564;
  assign n6566 = n6565 ^ n6338;
  assign n6687 = n6686 ^ n6566;
  assign n6556 = n2102 & n2448;
  assign n6557 = x89 & n2105;
  assign n6558 = x88 & n2112;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = x90 & n2381;
  assign n6561 = n6559 & ~n6560;
  assign n6562 = ~n6556 & n6561;
  assign n6563 = n6562 ^ x26;
  assign n6688 = n6687 ^ n6563;
  assign n6553 = n6434 ^ n6327;
  assign n6554 = ~n6435 & ~n6553;
  assign n6555 = n6554 ^ n6327;
  assign n6689 = n6688 ^ n6555;
  assign n6545 = n1746 & n2901;
  assign n6546 = x92 & n1750;
  assign n6547 = x91 & n1871;
  assign n6548 = ~n6546 & ~n6547;
  assign n6549 = x93 & n1873;
  assign n6550 = n6548 & ~n6549;
  assign n6551 = ~n6545 & n6550;
  assign n6552 = n6551 ^ x23;
  assign n6690 = n6689 ^ n6552;
  assign n6542 = n6436 ^ n6316;
  assign n6543 = n6437 & n6542;
  assign n6544 = n6543 ^ n6316;
  assign n6691 = n6690 ^ n6544;
  assign n6534 = n1404 & n3403;
  assign n6535 = x94 & n1514;
  assign n6536 = x95 & n1408;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = x96 & n1517;
  assign n6539 = n6537 & ~n6538;
  assign n6540 = ~n6534 & n6539;
  assign n6541 = n6540 ^ x20;
  assign n6692 = n6691 ^ n6541;
  assign n6531 = n6438 ^ n6305;
  assign n6532 = ~n6439 & ~n6531;
  assign n6533 = n6532 ^ n6305;
  assign n6693 = n6692 ^ n6533;
  assign n6523 = n1098 & n3943;
  assign n6524 = x98 & n1102;
  assign n6525 = x97 & n1198;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = x99 & n1201;
  assign n6528 = n6526 & ~n6527;
  assign n6529 = ~n6523 & n6528;
  assign n6530 = n6529 ^ x17;
  assign n6694 = n6693 ^ n6530;
  assign n6520 = n6440 ^ n6294;
  assign n6521 = n6441 & n6520;
  assign n6522 = n6521 ^ n6294;
  assign n6695 = n6694 ^ n6522;
  assign n6512 = n821 & n4509;
  assign n6513 = x100 & n898;
  assign n6514 = x101 & n824;
  assign n6515 = ~n6513 & ~n6514;
  assign n6516 = x102 & n901;
  assign n6517 = n6515 & ~n6516;
  assign n6518 = ~n6512 & n6517;
  assign n6519 = n6518 ^ x14;
  assign n6696 = n6695 ^ n6519;
  assign n6509 = n6442 ^ n6283;
  assign n6510 = ~n6443 & ~n6509;
  assign n6511 = n6510 ^ n6283;
  assign n6697 = n6696 ^ n6511;
  assign n6501 = n596 & n5117;
  assign n6502 = x104 & n601;
  assign n6503 = x103 & n673;
  assign n6504 = ~n6502 & ~n6503;
  assign n6505 = x105 & n676;
  assign n6506 = n6504 & ~n6505;
  assign n6507 = ~n6501 & n6506;
  assign n6508 = n6507 ^ x11;
  assign n6698 = n6697 ^ n6508;
  assign n6498 = n6444 ^ n6272;
  assign n6499 = n6445 & n6498;
  assign n6500 = n6499 ^ n6272;
  assign n6699 = n6698 ^ n6500;
  assign n6490 = n399 & n5792;
  assign n6491 = x106 & n478;
  assign n6492 = x108 & n470;
  assign n6493 = ~n6491 & ~n6492;
  assign n6494 = x107 & n402;
  assign n6495 = n6493 & ~n6494;
  assign n6496 = ~n6490 & n6495;
  assign n6497 = n6496 ^ x8;
  assign n6700 = n6699 ^ n6497;
  assign n6487 = n6446 ^ n6261;
  assign n6488 = ~n6447 & ~n6487;
  assign n6489 = n6488 ^ n6261;
  assign n6701 = n6700 ^ n6489;
  assign n6478 = n5782 ^ x111;
  assign n6479 = n239 & n6478;
  assign n6480 = x109 & n249;
  assign n6481 = x110 & n242;
  assign n6482 = ~n6480 & ~n6481;
  assign n6483 = x111 & n280;
  assign n6484 = n6482 & ~n6483;
  assign n6485 = ~n6479 & n6484;
  assign n6486 = n6485 ^ x5;
  assign n6702 = n6701 ^ n6486;
  assign n6475 = n6448 ^ n6248;
  assign n6476 = n6449 & ~n6475;
  assign n6477 = n6476 ^ n6248;
  assign n6703 = n6702 ^ n6477;
  assign n6464 = ~x112 & ~n6007;
  assign n6465 = x113 & ~n6464;
  assign n6466 = x112 & ~n6006;
  assign n6467 = ~x113 & ~n6466;
  assign n6468 = ~n6465 & ~n6467;
  assign n6469 = n169 & ~n6468;
  assign n6470 = n6469 ^ x1;
  assign n6471 = n6470 ^ x114;
  assign n6456 = x113 ^ x2;
  assign n6457 = n6456 ^ x112;
  assign n6458 = n6457 ^ n6456;
  assign n6459 = n6456 ^ x113;
  assign n6460 = ~n6458 & n6459;
  assign n6461 = n6460 ^ n6456;
  assign n6462 = ~x1 & n6461;
  assign n6463 = n6462 ^ n6456;
  assign n6472 = n6471 ^ n6463;
  assign n6473 = ~x0 & n6472;
  assign n6474 = n6473 ^ n6471;
  assign n6704 = n6703 ^ n6474;
  assign n6453 = n6450 ^ n6229;
  assign n6454 = ~n6451 & n6453;
  assign n6455 = n6454 ^ n6229;
  assign n6705 = n6704 ^ n6455;
  assign n6912 = n1149 & n4040;
  assign n6913 = x77 & n4267;
  assign n6914 = x78 & n4044;
  assign n6915 = ~n6913 & ~n6914;
  assign n6916 = x79 & n4270;
  assign n6917 = n6915 & ~n6916;
  assign n6918 = ~n6912 & n6917;
  assign n6919 = n6918 ^ x38;
  assign n6909 = n6679 ^ n6599;
  assign n6910 = ~n6680 & ~n6909;
  assign n6911 = n6910 ^ n6599;
  assign n6920 = n6919 ^ n6911;
  assign n6895 = n458 & n5942;
  assign n6896 = x69 & n5947;
  assign n6897 = x68 & n6186;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = x70 & n6406;
  assign n6900 = n6898 & ~n6899;
  assign n6901 = ~n6895 & n6900;
  assign n6902 = n6901 ^ x47;
  assign n6880 = n6411 ^ x50;
  assign n6881 = n6880 ^ n6411;
  assign n6882 = n6628 & n6881;
  assign n6883 = n6882 ^ n6411;
  assign n6884 = n6625 & n6883;
  assign n6885 = x65 & n6884;
  assign n6886 = x66 & n6630;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888 = n6191 & ~n6625;
  assign n6889 = x67 & n6888;
  assign n6890 = n6887 & ~n6889;
  assign n6891 = n285 & n6626;
  assign n6892 = n6890 & ~n6891;
  assign n6893 = n6892 ^ x50;
  assign n6878 = x51 ^ x50;
  assign n6879 = x64 & n6878;
  assign n6894 = n6893 ^ n6879;
  assign n6903 = n6902 ^ n6894;
  assign n6869 = n6621 & ~n6661;
  assign n6874 = n6643 & n6653;
  assign n6870 = n6664 ^ n6643;
  assign n6871 = n6653 ^ n6643;
  assign n6872 = n6870 & n6871;
  assign n6873 = n6872 ^ n6643;
  assign n6875 = n6874 ^ n6873;
  assign n6876 = ~n6869 & ~n6875;
  assign n6877 = n6876 ^ n6874;
  assign n6904 = n6903 ^ n6877;
  assign n6861 = ~n653 & n5262;
  assign n6862 = x72 & n5266;
  assign n6863 = x71 & n5488;
  assign n6864 = ~n6862 & ~n6863;
  assign n6865 = x73 & n5491;
  assign n6866 = n6864 & ~n6865;
  assign n6867 = ~n6861 & n6866;
  assign n6868 = n6867 ^ x44;
  assign n6905 = n6904 ^ n6868;
  assign n6858 = n6664 ^ n6615;
  assign n6859 = ~n6665 & ~n6858;
  assign n6860 = n6859 ^ n6618;
  assign n6906 = n6905 ^ n6860;
  assign n6850 = n870 & n4643;
  assign n6851 = x74 & n4653;
  assign n6852 = x75 & n4646;
  assign n6853 = ~n6851 & ~n6852;
  assign n6854 = x76 & n5046;
  assign n6855 = n6853 & ~n6854;
  assign n6856 = ~n6850 & n6855;
  assign n6857 = n6856 ^ x41;
  assign n6907 = n6906 ^ n6857;
  assign n6847 = n6677 ^ n6666;
  assign n6848 = ~n6678 & n6847;
  assign n6849 = n6848 ^ n6669;
  assign n6908 = n6907 ^ n6849;
  assign n6921 = n6920 ^ n6908;
  assign n6839 = n1454 & n3522;
  assign n6840 = x80 & n3699;
  assign n6841 = x82 & n3701;
  assign n6842 = ~n6840 & ~n6841;
  assign n6843 = x81 & n3526;
  assign n6844 = n6842 & ~n6843;
  assign n6845 = ~n6839 & n6844;
  assign n6846 = n6845 ^ x35;
  assign n6922 = n6921 ^ n6846;
  assign n6836 = n6681 ^ n6588;
  assign n6837 = n6682 & n6836;
  assign n6838 = n6837 ^ n6588;
  assign n6923 = n6922 ^ n6838;
  assign n6828 = n1801 & n3009;
  assign n6829 = x83 & n3181;
  assign n6830 = x84 & n3013;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = x85 & n3183;
  assign n6833 = n6831 & ~n6832;
  assign n6834 = ~n6828 & n6833;
  assign n6835 = n6834 ^ x32;
  assign n6924 = n6923 ^ n6835;
  assign n6825 = n6585 ^ n6577;
  assign n6826 = n6684 & n6825;
  assign n6827 = n6826 ^ n6683;
  assign n6925 = n6924 ^ n6827;
  assign n6817 = n2176 & n2527;
  assign n6818 = x86 & n2690;
  assign n6819 = x87 & n2530;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = x88 & n2693;
  assign n6822 = n6820 & ~n6821;
  assign n6823 = ~n6817 & n6822;
  assign n6824 = n6823 ^ x29;
  assign n6926 = n6925 ^ n6824;
  assign n6814 = n6685 ^ n6566;
  assign n6815 = n6686 & n6814;
  assign n6816 = n6815 ^ n6566;
  assign n6927 = n6926 ^ n6816;
  assign n6806 = n2102 & n2607;
  assign n6807 = x89 & n2112;
  assign n6808 = x91 & n2381;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = x90 & n2105;
  assign n6811 = n6809 & ~n6810;
  assign n6812 = ~n6806 & n6811;
  assign n6813 = n6812 ^ x26;
  assign n6928 = n6927 ^ n6813;
  assign n6803 = n6687 ^ n6555;
  assign n6804 = ~n6688 & ~n6803;
  assign n6805 = n6804 ^ n6555;
  assign n6929 = n6928 ^ n6805;
  assign n6795 = n1746 & n3078;
  assign n6796 = x93 & n1750;
  assign n6797 = x92 & n1871;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = x94 & n1873;
  assign n6800 = n6798 & ~n6799;
  assign n6801 = ~n6795 & n6800;
  assign n6802 = n6801 ^ x23;
  assign n6930 = n6929 ^ n6802;
  assign n6792 = n6689 ^ n6544;
  assign n6793 = n6690 & n6792;
  assign n6794 = n6793 ^ n6544;
  assign n6931 = n6930 ^ n6794;
  assign n6784 = n1404 & n3585;
  assign n6785 = x96 & n1408;
  assign n6786 = x95 & n1514;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = x97 & n1517;
  assign n6789 = n6787 & ~n6788;
  assign n6790 = ~n6784 & n6789;
  assign n6791 = n6790 ^ x20;
  assign n6932 = n6931 ^ n6791;
  assign n6781 = n6691 ^ n6533;
  assign n6782 = ~n6692 & ~n6781;
  assign n6783 = n6782 ^ n6533;
  assign n6933 = n6932 ^ n6783;
  assign n6773 = n1098 & n4141;
  assign n6774 = x98 & n1198;
  assign n6775 = x99 & n1102;
  assign n6776 = ~n6774 & ~n6775;
  assign n6777 = x100 & n1201;
  assign n6778 = n6776 & ~n6777;
  assign n6779 = ~n6773 & n6778;
  assign n6780 = n6779 ^ x17;
  assign n6934 = n6933 ^ n6780;
  assign n6770 = n6693 ^ n6522;
  assign n6771 = n6694 & n6770;
  assign n6772 = n6771 ^ n6522;
  assign n6935 = n6934 ^ n6772;
  assign n6762 = n821 & n4718;
  assign n6763 = x101 & n898;
  assign n6764 = x102 & n824;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = x103 & n901;
  assign n6767 = n6765 & ~n6766;
  assign n6768 = ~n6762 & n6767;
  assign n6769 = n6768 ^ x14;
  assign n6936 = n6935 ^ n6769;
  assign n6759 = n6695 ^ n6511;
  assign n6760 = ~n6696 & ~n6759;
  assign n6761 = n6760 ^ n6511;
  assign n6937 = n6936 ^ n6761;
  assign n6751 = n596 & n5351;
  assign n6752 = x104 & n673;
  assign n6753 = x105 & n601;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = x106 & n676;
  assign n6756 = n6754 & ~n6755;
  assign n6757 = ~n6751 & n6756;
  assign n6758 = n6757 ^ x11;
  assign n6938 = n6937 ^ n6758;
  assign n6748 = n6697 ^ n6500;
  assign n6749 = n6698 & n6748;
  assign n6750 = n6749 ^ n6500;
  assign n6939 = n6938 ^ n6750;
  assign n6740 = n399 & n6026;
  assign n6741 = x107 & n478;
  assign n6742 = x108 & n402;
  assign n6743 = ~n6741 & ~n6742;
  assign n6744 = x109 & n470;
  assign n6745 = n6743 & ~n6744;
  assign n6746 = ~n6740 & n6745;
  assign n6747 = n6746 ^ x8;
  assign n6940 = n6939 ^ n6747;
  assign n6737 = n6699 ^ n6489;
  assign n6738 = ~n6700 & ~n6737;
  assign n6739 = n6738 ^ n6489;
  assign n6941 = n6940 ^ n6739;
  assign n6728 = n6008 ^ x112;
  assign n6729 = n239 & n6728;
  assign n6730 = x110 & n249;
  assign n6731 = x111 & n242;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = x112 & n280;
  assign n6734 = n6732 & ~n6733;
  assign n6735 = ~n6729 & n6734;
  assign n6736 = n6735 ^ x5;
  assign n6942 = n6941 ^ n6736;
  assign n6725 = n6701 ^ n6477;
  assign n6726 = n6702 & ~n6725;
  assign n6727 = n6726 ^ n6477;
  assign n6943 = n6942 ^ n6727;
  assign n6714 = x114 ^ x2;
  assign n6715 = n6714 ^ x113;
  assign n6716 = n6715 ^ n6714;
  assign n6717 = n6714 ^ x114;
  assign n6718 = ~n6716 & n6717;
  assign n6719 = n6718 ^ n6714;
  assign n6720 = ~x1 & n6719;
  assign n6721 = n6720 ^ n6714;
  assign n6709 = x114 ^ x113;
  assign n6710 = ~n6468 & n6709;
  assign n6711 = n169 & ~n6710;
  assign n6712 = n6711 ^ x1;
  assign n6713 = n6712 ^ x115;
  assign n6722 = n6721 ^ n6713;
  assign n6723 = ~x0 & n6722;
  assign n6724 = n6723 ^ n6713;
  assign n6944 = n6943 ^ n6724;
  assign n6706 = n6703 ^ n6455;
  assign n6707 = ~n6704 & n6706;
  assign n6708 = n6707 ^ n6455;
  assign n6945 = n6944 ^ n6708;
  assign n7157 = n956 & n4643;
  assign n7158 = x75 & n4653;
  assign n7159 = x76 & n4646;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = x77 & n5046;
  assign n7162 = n7160 & ~n7161;
  assign n7163 = ~n7157 & n7162;
  assign n7164 = n7163 ^ x41;
  assign n7154 = n6906 ^ n6849;
  assign n7155 = n6907 & n7154;
  assign n7156 = n7155 ^ n6849;
  assign n7165 = n7164 ^ n7156;
  assign n7144 = ~n6869 & ~n6873;
  assign n7145 = n6903 & n7144;
  assign n7124 = ~n6874 & ~n6894;
  assign n7146 = ~n6869 & ~n6894;
  assign n7147 = ~n6902 & ~n7146;
  assign n7148 = ~n7124 & ~n7147;
  assign n7149 = ~n7145 & ~n7148;
  assign n7136 = n517 & n5942;
  assign n7137 = x70 & n5947;
  assign n7138 = x69 & n6186;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = x71 & n6406;
  assign n7141 = n7139 & ~n7140;
  assign n7142 = ~n7136 & n7141;
  assign n7143 = n7142 ^ x47;
  assign n7150 = n7149 ^ n7143;
  assign n7130 = x50 & x51;
  assign n7131 = n7130 ^ x52;
  assign n7132 = ~x64 & n7131;
  assign n7126 = x65 ^ x51;
  assign n7127 = n6878 & ~n7126;
  assign n7128 = n7127 ^ x50;
  assign n7129 = n7128 ^ x52;
  assign n7133 = n7132 ^ n7129;
  assign n7125 = ~n6893 & ~n7124;
  assign n7134 = n7133 ^ n7125;
  assign n7116 = n321 & n6626;
  assign n7117 = x67 & n6630;
  assign n7118 = x66 & n6884;
  assign n7119 = ~n7117 & ~n7118;
  assign n7120 = x68 & n6888;
  assign n7121 = n7119 & ~n7120;
  assign n7122 = ~n7116 & n7121;
  assign n7123 = n7122 ^ x50;
  assign n7135 = n7134 ^ n7123;
  assign n7151 = n7150 ^ n7135;
  assign n7108 = ~n721 & n5262;
  assign n7109 = x73 & n5266;
  assign n7110 = x72 & n5488;
  assign n7111 = ~n7109 & ~n7110;
  assign n7112 = x74 & n5491;
  assign n7113 = n7111 & ~n7112;
  assign n7114 = ~n7108 & n7113;
  assign n7115 = n7114 ^ x44;
  assign n7152 = n7151 ^ n7115;
  assign n7105 = n6904 ^ n6860;
  assign n7106 = ~n6905 & ~n7105;
  assign n7107 = n7106 ^ n6860;
  assign n7153 = n7152 ^ n7107;
  assign n7166 = n7165 ^ n7153;
  assign n7097 = n1242 & n4040;
  assign n7098 = x78 & n4267;
  assign n7099 = x80 & n4270;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = x79 & n4044;
  assign n7102 = n7100 & ~n7101;
  assign n7103 = ~n7097 & n7102;
  assign n7104 = n7103 ^ x38;
  assign n7167 = n7166 ^ n7104;
  assign n7094 = n6919 ^ n6908;
  assign n7095 = ~n6920 & ~n7094;
  assign n7096 = n7095 ^ n6911;
  assign n7168 = n7167 ^ n7096;
  assign n7086 = n1560 & n3522;
  assign n7087 = x81 & n3699;
  assign n7088 = x82 & n3526;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = x83 & n3701;
  assign n7091 = n7089 & ~n7090;
  assign n7092 = ~n7086 & n7091;
  assign n7093 = n7092 ^ x35;
  assign n7169 = n7168 ^ n7093;
  assign n7083 = n6921 ^ n6838;
  assign n7084 = n6922 & n7083;
  assign n7085 = n7084 ^ n6838;
  assign n7170 = n7169 ^ n7085;
  assign n7075 = n1920 & n3009;
  assign n7076 = x85 & n3013;
  assign n7077 = x84 & n3181;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = x86 & n3183;
  assign n7080 = n7078 & ~n7079;
  assign n7081 = ~n7075 & n7080;
  assign n7082 = n7081 ^ x32;
  assign n7171 = n7170 ^ n7082;
  assign n7072 = n6835 ^ n6827;
  assign n7073 = n6924 & ~n7072;
  assign n7074 = n7073 ^ n6923;
  assign n7172 = n7171 ^ n7074;
  assign n7064 = n2310 & n2527;
  assign n7065 = x88 & n2530;
  assign n7066 = x87 & n2690;
  assign n7067 = ~n7065 & ~n7066;
  assign n7068 = x89 & n2693;
  assign n7069 = n7067 & ~n7068;
  assign n7070 = ~n7064 & n7069;
  assign n7071 = n7070 ^ x29;
  assign n7173 = n7172 ^ n7071;
  assign n7061 = n6925 ^ n6816;
  assign n7062 = ~n6926 & ~n7061;
  assign n7063 = n7062 ^ n6816;
  assign n7174 = n7173 ^ n7063;
  assign n7053 = n2102 & n2755;
  assign n7054 = x90 & n2112;
  assign n7055 = x92 & n2381;
  assign n7056 = ~n7054 & ~n7055;
  assign n7057 = x91 & n2105;
  assign n7058 = n7056 & ~n7057;
  assign n7059 = ~n7053 & n7058;
  assign n7060 = n7059 ^ x26;
  assign n7175 = n7174 ^ n7060;
  assign n7050 = n6927 ^ n6805;
  assign n7051 = n6928 & n7050;
  assign n7052 = n7051 ^ n6805;
  assign n7176 = n7175 ^ n7052;
  assign n7042 = n1746 & n3247;
  assign n7043 = x94 & n1750;
  assign n7044 = x93 & n1871;
  assign n7045 = ~n7043 & ~n7044;
  assign n7046 = x95 & n1873;
  assign n7047 = n7045 & ~n7046;
  assign n7048 = ~n7042 & n7047;
  assign n7049 = n7048 ^ x23;
  assign n7177 = n7176 ^ n7049;
  assign n7039 = n6929 ^ n6794;
  assign n7040 = ~n6930 & ~n7039;
  assign n7041 = n7040 ^ n6794;
  assign n7178 = n7177 ^ n7041;
  assign n7031 = n1404 & n3763;
  assign n7032 = x96 & n1514;
  assign n7033 = x98 & n1517;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = x97 & n1408;
  assign n7036 = n7034 & ~n7035;
  assign n7037 = ~n7031 & n7036;
  assign n7038 = n7037 ^ x20;
  assign n7179 = n7178 ^ n7038;
  assign n7028 = n6931 ^ n6783;
  assign n7029 = n6932 & n7028;
  assign n7030 = n7029 ^ n6783;
  assign n7180 = n7179 ^ n7030;
  assign n7020 = n1098 & n4323;
  assign n7021 = x100 & n1102;
  assign n7022 = x99 & n1198;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = x101 & n1201;
  assign n7025 = n7023 & ~n7024;
  assign n7026 = ~n7020 & n7025;
  assign n7027 = n7026 ^ x17;
  assign n7181 = n7180 ^ n7027;
  assign n7017 = n6933 ^ n6772;
  assign n7018 = ~n6934 & ~n7017;
  assign n7019 = n7018 ^ n6772;
  assign n7182 = n7181 ^ n7019;
  assign n7009 = n821 & n4912;
  assign n7010 = x103 & n824;
  assign n7011 = x102 & n898;
  assign n7012 = ~n7010 & ~n7011;
  assign n7013 = x104 & n901;
  assign n7014 = n7012 & ~n7013;
  assign n7015 = ~n7009 & n7014;
  assign n7016 = n7015 ^ x14;
  assign n7183 = n7182 ^ n7016;
  assign n7006 = n6935 ^ n6761;
  assign n7007 = n6936 & n7006;
  assign n7008 = n7007 ^ n6761;
  assign n7184 = n7183 ^ n7008;
  assign n6998 = n596 & n5578;
  assign n6999 = x105 & n673;
  assign n7000 = x106 & n601;
  assign n7001 = ~n6999 & ~n7000;
  assign n7002 = x107 & n676;
  assign n7003 = n7001 & ~n7002;
  assign n7004 = ~n6998 & n7003;
  assign n7005 = n7004 ^ x11;
  assign n7185 = n7184 ^ n7005;
  assign n6995 = n6937 ^ n6750;
  assign n6996 = ~n6938 & ~n6995;
  assign n6997 = n6996 ^ n6750;
  assign n7186 = n7185 ^ n6997;
  assign n6987 = n399 & n6250;
  assign n6988 = x108 & n478;
  assign n6989 = x109 & n402;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = x110 & n470;
  assign n6992 = n6990 & ~n6991;
  assign n6993 = ~n6987 & n6992;
  assign n6994 = n6993 ^ x8;
  assign n7187 = n7186 ^ n6994;
  assign n6984 = n6939 ^ n6739;
  assign n6985 = n6940 & n6984;
  assign n6986 = n6985 ^ n6739;
  assign n7188 = n7187 ^ n6986;
  assign n6975 = n6233 ^ x113;
  assign n6976 = n239 & n6975;
  assign n6977 = x111 & n249;
  assign n6978 = x112 & n242;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = x113 & n280;
  assign n6981 = n6979 & ~n6980;
  assign n6982 = ~n6976 & n6981;
  assign n6983 = n6982 ^ x5;
  assign n7189 = n7188 ^ n6983;
  assign n6972 = n6941 ^ n6727;
  assign n6973 = ~n6942 & n6972;
  assign n6974 = n6973 ^ n6727;
  assign n7190 = n7189 ^ n6974;
  assign n6961 = ~x114 & ~n6465;
  assign n6962 = x115 & ~n6961;
  assign n6963 = x114 & ~n6467;
  assign n6964 = ~x115 & ~n6963;
  assign n6965 = ~n6962 & ~n6964;
  assign n6966 = n169 & ~n6965;
  assign n6967 = n6966 ^ x1;
  assign n6968 = n6967 ^ x116;
  assign n6949 = x115 ^ x2;
  assign n6950 = n6949 ^ x1;
  assign n6951 = n6950 ^ n6949;
  assign n6952 = n6951 ^ x0;
  assign n6953 = n6949 ^ x115;
  assign n6954 = n6953 ^ x114;
  assign n6955 = ~x114 & ~n6954;
  assign n6956 = n6955 ^ n6949;
  assign n6957 = n6956 ^ x114;
  assign n6958 = n6952 & ~n6957;
  assign n6959 = n6958 ^ n6955;
  assign n6960 = n6959 ^ x114;
  assign n6969 = n6968 ^ n6960;
  assign n6970 = ~x0 & ~n6969;
  assign n6971 = n6970 ^ n6968;
  assign n7191 = n7190 ^ n6971;
  assign n6946 = n6943 ^ n6708;
  assign n6947 = n6944 & ~n6946;
  assign n6948 = n6947 ^ n6708;
  assign n7192 = n7191 ^ n6948;
  assign n7417 = x52 ^ x50;
  assign n7418 = x64 & n7417;
  assign n7419 = n7418 ^ n233;
  assign n7420 = ~n6878 & ~n7419;
  assign n7421 = n7420 ^ n233;
  assign n7422 = x53 & n7421;
  assign n7394 = x53 ^ x52;
  assign n7395 = n6878 & n7394;
  assign n7396 = n142 & n7395;
  assign n7397 = ~x50 & ~x51;
  assign n7398 = n7397 ^ n7130;
  assign n7399 = x52 & n7398;
  assign n7400 = n7399 ^ n7130;
  assign n7401 = ~n7396 & ~n7400;
  assign n7402 = x65 & ~n7401;
  assign n7403 = n152 & n7394;
  assign n7404 = x66 & n6878;
  assign n7405 = ~n7403 & n7404;
  assign n7406 = ~n7402 & ~n7405;
  assign n7407 = n7406 ^ x53;
  assign n7411 = x52 & ~x53;
  assign n7412 = n7130 & n7411;
  assign n7413 = x64 & n7412;
  assign n7408 = ~x52 & x64;
  assign n7409 = n7397 & n7408;
  assign n7410 = x53 & n7409;
  assign n7414 = n7413 ^ n7410;
  assign n7415 = ~n7407 & ~n7414;
  assign n7416 = n7415 ^ n7413;
  assign n7423 = n7422 ^ n7416;
  assign n7386 = n420 & n6626;
  assign n7387 = x68 & n6630;
  assign n7388 = x67 & n6884;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = x69 & n6888;
  assign n7391 = n7389 & ~n7390;
  assign n7392 = ~n7386 & n7391;
  assign n7393 = n7392 ^ x50;
  assign n7424 = n7423 ^ n7393;
  assign n7383 = n7133 ^ n7123;
  assign n7384 = n7134 & n7383;
  assign n7385 = n7384 ^ n7125;
  assign n7425 = n7424 ^ n7385;
  assign n7375 = n575 & n5942;
  assign n7376 = x71 & n5947;
  assign n7377 = x70 & n6186;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = x72 & n6406;
  assign n7380 = n7378 & ~n7379;
  assign n7381 = ~n7375 & n7380;
  assign n7382 = n7381 ^ x47;
  assign n7426 = n7425 ^ n7382;
  assign n7372 = n7143 ^ n7135;
  assign n7373 = ~n7150 & ~n7372;
  assign n7374 = n7373 ^ n7149;
  assign n7427 = n7426 ^ n7374;
  assign n7364 = n789 & n5262;
  assign n7365 = x74 & n5266;
  assign n7366 = x75 & n5491;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = x73 & n5488;
  assign n7369 = n7367 & ~n7368;
  assign n7370 = ~n7364 & n7369;
  assign n7371 = n7370 ^ x44;
  assign n7428 = n7427 ^ n7371;
  assign n7361 = n7151 ^ n7107;
  assign n7362 = n7152 & n7361;
  assign n7363 = n7362 ^ n7107;
  assign n7429 = n7428 ^ n7363;
  assign n7353 = n1041 & n4643;
  assign n7354 = x76 & n4653;
  assign n7355 = x78 & n5046;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = x77 & n4646;
  assign n7358 = n7356 & ~n7357;
  assign n7359 = ~n7353 & n7358;
  assign n7360 = n7359 ^ x41;
  assign n7430 = n7429 ^ n7360;
  assign n7350 = n7164 ^ n7153;
  assign n7351 = ~n7165 & ~n7350;
  assign n7352 = n7351 ^ n7156;
  assign n7431 = n7430 ^ n7352;
  assign n7347 = n7166 ^ n7096;
  assign n7348 = n7167 & n7347;
  assign n7349 = n7348 ^ n7096;
  assign n7432 = n7431 ^ n7349;
  assign n7339 = n1340 & n4040;
  assign n7340 = x80 & n4044;
  assign n7341 = x81 & n4270;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = x79 & n4267;
  assign n7344 = n7342 & ~n7343;
  assign n7345 = ~n7339 & n7344;
  assign n7346 = n7345 ^ x38;
  assign n7433 = n7432 ^ n7346;
  assign n7331 = n1667 & n3522;
  assign n7332 = x82 & n3699;
  assign n7333 = x83 & n3526;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = x84 & n3701;
  assign n7336 = n7334 & ~n7335;
  assign n7337 = ~n7331 & n7336;
  assign n7338 = n7337 ^ x35;
  assign n7434 = n7433 ^ n7338;
  assign n7328 = n7168 ^ n7085;
  assign n7329 = ~n7169 & ~n7328;
  assign n7330 = n7329 ^ n7085;
  assign n7435 = n7434 ^ n7330;
  assign n7320 = n2039 & n3009;
  assign n7321 = x86 & n3013;
  assign n7322 = x85 & n3181;
  assign n7323 = ~n7321 & ~n7322;
  assign n7324 = x87 & n3183;
  assign n7325 = n7323 & ~n7324;
  assign n7326 = ~n7320 & n7325;
  assign n7327 = n7326 ^ x32;
  assign n7436 = n7435 ^ n7327;
  assign n7317 = n7082 ^ n7074;
  assign n7318 = ~n7171 & ~n7317;
  assign n7319 = n7318 ^ n7170;
  assign n7437 = n7436 ^ n7319;
  assign n7309 = n2448 & n2527;
  assign n7310 = x88 & n2690;
  assign n7311 = x90 & n2693;
  assign n7312 = ~n7310 & ~n7311;
  assign n7313 = x89 & n2530;
  assign n7314 = n7312 & ~n7313;
  assign n7315 = ~n7309 & n7314;
  assign n7316 = n7315 ^ x29;
  assign n7438 = n7437 ^ n7316;
  assign n7306 = n7172 ^ n7063;
  assign n7307 = n7173 & n7306;
  assign n7308 = n7307 ^ n7063;
  assign n7439 = n7438 ^ n7308;
  assign n7298 = n2102 & n2901;
  assign n7299 = x91 & n2112;
  assign n7300 = x93 & n2381;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = x92 & n2105;
  assign n7303 = n7301 & ~n7302;
  assign n7304 = ~n7298 & n7303;
  assign n7305 = n7304 ^ x26;
  assign n7440 = n7439 ^ n7305;
  assign n7295 = n7174 ^ n7052;
  assign n7296 = ~n7175 & ~n7295;
  assign n7297 = n7296 ^ n7052;
  assign n7441 = n7440 ^ n7297;
  assign n7287 = n1746 & n3403;
  assign n7288 = x94 & n1871;
  assign n7289 = x95 & n1750;
  assign n7290 = ~n7288 & ~n7289;
  assign n7291 = x96 & n1873;
  assign n7292 = n7290 & ~n7291;
  assign n7293 = ~n7287 & n7292;
  assign n7294 = n7293 ^ x23;
  assign n7442 = n7441 ^ n7294;
  assign n7284 = n7176 ^ n7041;
  assign n7285 = n7177 & n7284;
  assign n7286 = n7285 ^ n7041;
  assign n7443 = n7442 ^ n7286;
  assign n7276 = n1404 & n3943;
  assign n7277 = x98 & n1408;
  assign n7278 = x97 & n1514;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = x99 & n1517;
  assign n7281 = n7279 & ~n7280;
  assign n7282 = ~n7276 & n7281;
  assign n7283 = n7282 ^ x20;
  assign n7444 = n7443 ^ n7283;
  assign n7273 = n7178 ^ n7030;
  assign n7274 = ~n7179 & ~n7273;
  assign n7275 = n7274 ^ n7030;
  assign n7445 = n7444 ^ n7275;
  assign n7265 = n1098 & n4509;
  assign n7266 = x101 & n1102;
  assign n7267 = x100 & n1198;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = x102 & n1201;
  assign n7270 = n7268 & ~n7269;
  assign n7271 = ~n7265 & n7270;
  assign n7272 = n7271 ^ x17;
  assign n7446 = n7445 ^ n7272;
  assign n7262 = n7180 ^ n7019;
  assign n7263 = n7181 & n7262;
  assign n7264 = n7263 ^ n7019;
  assign n7447 = n7446 ^ n7264;
  assign n7254 = n821 & n5117;
  assign n7255 = x103 & n898;
  assign n7256 = x105 & n901;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = x104 & n824;
  assign n7259 = n7257 & ~n7258;
  assign n7260 = ~n7254 & n7259;
  assign n7261 = n7260 ^ x14;
  assign n7448 = n7447 ^ n7261;
  assign n7251 = n7182 ^ n7008;
  assign n7252 = ~n7183 & ~n7251;
  assign n7253 = n7252 ^ n7008;
  assign n7449 = n7448 ^ n7253;
  assign n7243 = n596 & n5792;
  assign n7244 = x106 & n673;
  assign n7245 = x107 & n601;
  assign n7246 = ~n7244 & ~n7245;
  assign n7247 = x108 & n676;
  assign n7248 = n7246 & ~n7247;
  assign n7249 = ~n7243 & n7248;
  assign n7250 = n7249 ^ x11;
  assign n7450 = n7449 ^ n7250;
  assign n7240 = n7184 ^ n6997;
  assign n7241 = n7185 & n7240;
  assign n7242 = n7241 ^ n6997;
  assign n7451 = n7450 ^ n7242;
  assign n7232 = n399 & n6478;
  assign n7233 = x109 & n478;
  assign n7234 = x111 & n470;
  assign n7235 = ~n7233 & ~n7234;
  assign n7236 = x110 & n402;
  assign n7237 = n7235 & ~n7236;
  assign n7238 = ~n7232 & n7237;
  assign n7239 = n7238 ^ x8;
  assign n7452 = n7451 ^ n7239;
  assign n7229 = n7186 ^ n6986;
  assign n7230 = ~n7187 & ~n7229;
  assign n7231 = n7230 ^ n6986;
  assign n7453 = n7452 ^ n7231;
  assign n7220 = n6468 ^ x114;
  assign n7221 = n239 & n7220;
  assign n7222 = x112 & n249;
  assign n7223 = x114 & n280;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = x113 & n242;
  assign n7226 = n7224 & ~n7225;
  assign n7227 = ~n7221 & n7226;
  assign n7228 = n7227 ^ x5;
  assign n7454 = n7453 ^ n7228;
  assign n7217 = n7188 ^ n6974;
  assign n7218 = n7189 & ~n7217;
  assign n7219 = n7218 ^ n6974;
  assign n7455 = n7454 ^ n7219;
  assign n7208 = ~x116 & ~n6962;
  assign n7209 = x116 & ~n6964;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = n169 & ~n7210;
  assign n7212 = n7211 ^ x1;
  assign n7213 = n7212 ^ x117;
  assign n7196 = x116 ^ x2;
  assign n7197 = n7196 ^ x1;
  assign n7198 = n7197 ^ n7196;
  assign n7199 = n7198 ^ x0;
  assign n7200 = n7196 ^ x116;
  assign n7201 = n7200 ^ x115;
  assign n7202 = ~x115 & ~n7201;
  assign n7203 = n7202 ^ n7196;
  assign n7204 = n7203 ^ x115;
  assign n7205 = n7199 & ~n7204;
  assign n7206 = n7205 ^ n7202;
  assign n7207 = n7206 ^ x115;
  assign n7214 = n7213 ^ n7207;
  assign n7215 = ~x0 & ~n7214;
  assign n7216 = n7215 ^ n7213;
  assign n7456 = n7455 ^ n7216;
  assign n7193 = n7190 ^ n6948;
  assign n7194 = ~n7191 & n7193;
  assign n7195 = n7194 ^ n6948;
  assign n7457 = n7456 ^ n7195;
  assign n7672 = n1149 & n4643;
  assign n7673 = x77 & n4653;
  assign n7674 = x79 & n5046;
  assign n7675 = ~n7673 & ~n7674;
  assign n7676 = x78 & n4646;
  assign n7677 = n7675 & ~n7676;
  assign n7678 = ~n7672 & n7677;
  assign n7679 = n7678 ^ x41;
  assign n7669 = n7429 ^ n7352;
  assign n7670 = ~n7430 & ~n7669;
  assign n7671 = n7670 ^ n7352;
  assign n7680 = n7679 ^ n7671;
  assign n7661 = n7416 & n7422;
  assign n7646 = n7130 ^ x53;
  assign n7647 = n7646 ^ n7130;
  assign n7648 = n7398 & n7647;
  assign n7649 = n7648 ^ n7130;
  assign n7650 = n7394 & n7649;
  assign n7651 = x65 & n7650;
  assign n7652 = n6878 & ~n7394;
  assign n7653 = x67 & n7652;
  assign n7654 = ~n7651 & ~n7653;
  assign n7655 = x66 & n7400;
  assign n7656 = n7654 & ~n7655;
  assign n7657 = n285 & n7395;
  assign n7658 = n7656 & ~n7657;
  assign n7659 = n7658 ^ x53;
  assign n7644 = x54 ^ x53;
  assign n7645 = x64 & n7644;
  assign n7660 = n7659 ^ n7645;
  assign n7662 = n7661 ^ n7660;
  assign n7636 = n458 & n6626;
  assign n7637 = x68 & n6884;
  assign n7638 = x69 & n6630;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = x70 & n6888;
  assign n7641 = n7639 & ~n7640;
  assign n7642 = ~n7636 & n7641;
  assign n7643 = n7642 ^ x50;
  assign n7663 = n7662 ^ n7643;
  assign n7633 = n7423 ^ n7385;
  assign n7634 = n7424 & n7633;
  assign n7635 = n7634 ^ n7385;
  assign n7664 = n7663 ^ n7635;
  assign n7625 = ~n653 & n5942;
  assign n7626 = x72 & n5947;
  assign n7627 = x71 & n6186;
  assign n7628 = ~n7626 & ~n7627;
  assign n7629 = x73 & n6406;
  assign n7630 = n7628 & ~n7629;
  assign n7631 = ~n7625 & n7630;
  assign n7632 = n7631 ^ x47;
  assign n7665 = n7664 ^ n7632;
  assign n7622 = n7425 ^ n7374;
  assign n7623 = ~n7426 & ~n7622;
  assign n7624 = n7623 ^ n7374;
  assign n7666 = n7665 ^ n7624;
  assign n7614 = n870 & n5262;
  assign n7615 = x74 & n5488;
  assign n7616 = x75 & n5266;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = x76 & n5491;
  assign n7619 = n7617 & ~n7618;
  assign n7620 = ~n7614 & n7619;
  assign n7621 = n7620 ^ x44;
  assign n7667 = n7666 ^ n7621;
  assign n7611 = n7427 ^ n7363;
  assign n7612 = n7428 & n7611;
  assign n7613 = n7612 ^ n7363;
  assign n7668 = n7667 ^ n7613;
  assign n7681 = n7680 ^ n7668;
  assign n7603 = n1454 & n4040;
  assign n7604 = x80 & n4267;
  assign n7605 = x82 & n4270;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = x81 & n4044;
  assign n7608 = n7606 & ~n7607;
  assign n7609 = ~n7603 & n7608;
  assign n7610 = n7609 ^ x38;
  assign n7682 = n7681 ^ n7610;
  assign n7600 = n7431 ^ n7346;
  assign n7601 = n7432 & n7600;
  assign n7602 = n7601 ^ n7349;
  assign n7683 = n7682 ^ n7602;
  assign n7592 = n1801 & n3522;
  assign n7593 = x83 & n3699;
  assign n7594 = x85 & n3701;
  assign n7595 = ~n7593 & ~n7594;
  assign n7596 = x84 & n3526;
  assign n7597 = n7595 & ~n7596;
  assign n7598 = ~n7592 & n7597;
  assign n7599 = n7598 ^ x35;
  assign n7684 = n7683 ^ n7599;
  assign n7589 = n7433 ^ n7330;
  assign n7590 = ~n7434 & ~n7589;
  assign n7591 = n7590 ^ n7330;
  assign n7685 = n7684 ^ n7591;
  assign n7581 = n2176 & n3009;
  assign n7582 = x87 & n3013;
  assign n7583 = x86 & n3181;
  assign n7584 = ~n7582 & ~n7583;
  assign n7585 = x88 & n3183;
  assign n7586 = n7584 & ~n7585;
  assign n7587 = ~n7581 & n7586;
  assign n7588 = n7587 ^ x32;
  assign n7686 = n7685 ^ n7588;
  assign n7578 = n7435 ^ n7319;
  assign n7579 = n7436 & n7578;
  assign n7580 = n7579 ^ n7319;
  assign n7687 = n7686 ^ n7580;
  assign n7570 = n2527 & n2607;
  assign n7571 = x89 & n2690;
  assign n7572 = x90 & n2530;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = x91 & n2693;
  assign n7575 = n7573 & ~n7574;
  assign n7576 = ~n7570 & n7575;
  assign n7577 = n7576 ^ x29;
  assign n7688 = n7687 ^ n7577;
  assign n7567 = n7437 ^ n7308;
  assign n7568 = ~n7438 & ~n7567;
  assign n7569 = n7568 ^ n7308;
  assign n7689 = n7688 ^ n7569;
  assign n7559 = n2102 & n3078;
  assign n7560 = x93 & n2105;
  assign n7561 = x92 & n2112;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = x94 & n2381;
  assign n7564 = n7562 & ~n7563;
  assign n7565 = ~n7559 & n7564;
  assign n7566 = n7565 ^ x26;
  assign n7690 = n7689 ^ n7566;
  assign n7556 = n7439 ^ n7297;
  assign n7557 = n7440 & n7556;
  assign n7558 = n7557 ^ n7297;
  assign n7691 = n7690 ^ n7558;
  assign n7548 = n1746 & n3585;
  assign n7549 = x96 & n1750;
  assign n7550 = x95 & n1871;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = x97 & n1873;
  assign n7553 = n7551 & ~n7552;
  assign n7554 = ~n7548 & n7553;
  assign n7555 = n7554 ^ x23;
  assign n7692 = n7691 ^ n7555;
  assign n7545 = n7441 ^ n7286;
  assign n7546 = ~n7442 & ~n7545;
  assign n7547 = n7546 ^ n7286;
  assign n7693 = n7692 ^ n7547;
  assign n7537 = n1404 & n4141;
  assign n7538 = x98 & n1514;
  assign n7539 = x99 & n1408;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = x100 & n1517;
  assign n7542 = n7540 & ~n7541;
  assign n7543 = ~n7537 & n7542;
  assign n7544 = n7543 ^ x20;
  assign n7694 = n7693 ^ n7544;
  assign n7534 = n7443 ^ n7275;
  assign n7535 = n7444 & n7534;
  assign n7536 = n7535 ^ n7275;
  assign n7695 = n7694 ^ n7536;
  assign n7526 = n1098 & n4718;
  assign n7527 = x102 & n1102;
  assign n7528 = x101 & n1198;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = x103 & n1201;
  assign n7531 = n7529 & ~n7530;
  assign n7532 = ~n7526 & n7531;
  assign n7533 = n7532 ^ x17;
  assign n7696 = n7695 ^ n7533;
  assign n7523 = n7445 ^ n7264;
  assign n7524 = ~n7446 & ~n7523;
  assign n7525 = n7524 ^ n7264;
  assign n7697 = n7696 ^ n7525;
  assign n7515 = n821 & n5351;
  assign n7516 = x104 & n898;
  assign n7517 = x106 & n901;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = x105 & n824;
  assign n7520 = n7518 & ~n7519;
  assign n7521 = ~n7515 & n7520;
  assign n7522 = n7521 ^ x14;
  assign n7698 = n7697 ^ n7522;
  assign n7507 = n596 & n6026;
  assign n7508 = x107 & n673;
  assign n7509 = x108 & n601;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = x109 & n676;
  assign n7512 = n7510 & ~n7511;
  assign n7513 = ~n7507 & n7512;
  assign n7514 = n7513 ^ x11;
  assign n7699 = n7698 ^ n7514;
  assign n7504 = n7447 ^ n7253;
  assign n7505 = n7448 & n7504;
  assign n7506 = n7505 ^ n7253;
  assign n7700 = n7699 ^ n7506;
  assign n7501 = n7449 ^ n7242;
  assign n7502 = ~n7450 & ~n7501;
  assign n7503 = n7502 ^ n7242;
  assign n7701 = n7700 ^ n7503;
  assign n7493 = n399 & n6728;
  assign n7494 = x110 & n478;
  assign n7495 = x112 & n470;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = x111 & n402;
  assign n7498 = n7496 & ~n7497;
  assign n7499 = ~n7493 & n7498;
  assign n7500 = n7499 ^ x8;
  assign n7702 = n7701 ^ n7500;
  assign n7490 = n7451 ^ n7231;
  assign n7491 = n7452 & n7490;
  assign n7492 = n7491 ^ n7231;
  assign n7703 = n7702 ^ n7492;
  assign n7481 = n6710 ^ x115;
  assign n7482 = n239 & n7481;
  assign n7483 = x113 & n249;
  assign n7484 = x115 & n280;
  assign n7485 = ~n7483 & ~n7484;
  assign n7486 = x114 & n242;
  assign n7487 = n7485 & ~n7486;
  assign n7488 = ~n7482 & n7487;
  assign n7489 = n7488 ^ x5;
  assign n7704 = n7703 ^ n7489;
  assign n7478 = n7453 ^ n7219;
  assign n7479 = ~n7454 & n7478;
  assign n7480 = n7479 ^ n7219;
  assign n7705 = n7704 ^ n7480;
  assign n7462 = x117 & ~n7208;
  assign n7463 = ~x117 & ~n7209;
  assign n7464 = ~n7462 & ~n7463;
  assign n7465 = n169 & ~n7464;
  assign n7466 = n7465 ^ x1;
  assign n7467 = n7466 ^ x118;
  assign n7461 = ~x116 & n197;
  assign n7468 = n7467 ^ n7461;
  assign n7469 = n7468 ^ n7467;
  assign n7470 = x117 ^ x2;
  assign n7471 = x1 & n7470;
  assign n7472 = n7471 ^ n7467;
  assign n7473 = n7472 ^ n7467;
  assign n7474 = ~n7469 & ~n7473;
  assign n7475 = n7474 ^ n7467;
  assign n7476 = ~x0 & ~n7475;
  assign n7477 = n7476 ^ n7467;
  assign n7706 = n7705 ^ n7477;
  assign n7458 = n7455 ^ n7195;
  assign n7459 = n7456 & ~n7458;
  assign n7460 = n7459 ^ n7195;
  assign n7707 = n7706 ^ n7460;
  assign n7922 = n956 & n5262;
  assign n7923 = x75 & n5488;
  assign n7924 = x77 & n5491;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = x76 & n5266;
  assign n7927 = n7925 & ~n7926;
  assign n7928 = ~n7922 & n7927;
  assign n7929 = n7928 ^ x44;
  assign n7919 = n7666 ^ n7613;
  assign n7920 = ~n7667 & ~n7919;
  assign n7921 = n7920 ^ n7613;
  assign n7930 = n7929 ^ n7921;
  assign n7912 = ~n7645 & ~n7661;
  assign n7913 = ~n7659 & ~n7912;
  assign n7903 = n321 & n7395;
  assign n7904 = x67 & n7400;
  assign n7905 = x66 & n7650;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = x68 & n7652;
  assign n7908 = n7906 & ~n7907;
  assign n7909 = ~n7903 & n7908;
  assign n7910 = n7909 ^ x53;
  assign n7898 = x65 ^ x54;
  assign n7899 = n7644 & ~n7898;
  assign n7900 = n7899 ^ x53;
  assign n7901 = n7900 ^ x55;
  assign n7895 = x53 & x54;
  assign n7896 = n7895 ^ x55;
  assign n7897 = ~x64 & n7896;
  assign n7902 = n7901 ^ n7897;
  assign n7911 = n7910 ^ n7902;
  assign n7914 = n7913 ^ n7911;
  assign n7887 = n517 & n6626;
  assign n7888 = x70 & n6630;
  assign n7889 = x69 & n6884;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = x71 & n6888;
  assign n7892 = n7890 & ~n7891;
  assign n7893 = ~n7887 & n7892;
  assign n7894 = n7893 ^ x50;
  assign n7915 = n7914 ^ n7894;
  assign n7884 = n7662 ^ n7635;
  assign n7885 = ~n7663 & ~n7884;
  assign n7886 = n7885 ^ n7635;
  assign n7916 = n7915 ^ n7886;
  assign n7876 = ~n721 & n5942;
  assign n7877 = x73 & n5947;
  assign n7878 = x72 & n6186;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = x74 & n6406;
  assign n7881 = n7879 & ~n7880;
  assign n7882 = ~n7876 & n7881;
  assign n7883 = n7882 ^ x47;
  assign n7917 = n7916 ^ n7883;
  assign n7873 = n7664 ^ n7624;
  assign n7874 = n7665 & n7873;
  assign n7875 = n7874 ^ n7624;
  assign n7918 = n7917 ^ n7875;
  assign n7931 = n7930 ^ n7918;
  assign n7865 = n1242 & n4643;
  assign n7866 = x78 & n4653;
  assign n7867 = x79 & n4646;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = x80 & n5046;
  assign n7870 = n7868 & ~n7869;
  assign n7871 = ~n7865 & n7870;
  assign n7872 = n7871 ^ x41;
  assign n7932 = n7931 ^ n7872;
  assign n7862 = n7679 ^ n7668;
  assign n7863 = ~n7680 & n7862;
  assign n7864 = n7863 ^ n7671;
  assign n7933 = n7932 ^ n7864;
  assign n7854 = n1560 & n4040;
  assign n7855 = x81 & n4267;
  assign n7856 = x82 & n4044;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = x83 & n4270;
  assign n7859 = n7857 & ~n7858;
  assign n7860 = ~n7854 & n7859;
  assign n7861 = n7860 ^ x38;
  assign n7934 = n7933 ^ n7861;
  assign n7851 = n7681 ^ n7602;
  assign n7852 = ~n7682 & ~n7851;
  assign n7853 = n7852 ^ n7602;
  assign n7935 = n7934 ^ n7853;
  assign n7843 = n1920 & n3522;
  assign n7844 = x84 & n3699;
  assign n7845 = x86 & n3701;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = x85 & n3526;
  assign n7848 = n7846 & ~n7847;
  assign n7849 = ~n7843 & n7848;
  assign n7850 = n7849 ^ x35;
  assign n7936 = n7935 ^ n7850;
  assign n7840 = n7683 ^ n7591;
  assign n7841 = n7684 & n7840;
  assign n7842 = n7841 ^ n7591;
  assign n7937 = n7936 ^ n7842;
  assign n7832 = n2310 & n3009;
  assign n7833 = x87 & n3181;
  assign n7834 = x88 & n3013;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = x89 & n3183;
  assign n7837 = n7835 & ~n7836;
  assign n7838 = ~n7832 & n7837;
  assign n7839 = n7838 ^ x32;
  assign n7938 = n7937 ^ n7839;
  assign n7829 = n7685 ^ n7580;
  assign n7830 = ~n7686 & ~n7829;
  assign n7831 = n7830 ^ n7580;
  assign n7939 = n7938 ^ n7831;
  assign n7821 = n2527 & n2755;
  assign n7822 = x90 & n2690;
  assign n7823 = x91 & n2530;
  assign n7824 = ~n7822 & ~n7823;
  assign n7825 = x92 & n2693;
  assign n7826 = n7824 & ~n7825;
  assign n7827 = ~n7821 & n7826;
  assign n7828 = n7827 ^ x29;
  assign n7940 = n7939 ^ n7828;
  assign n7818 = n7687 ^ n7569;
  assign n7819 = n7688 & n7818;
  assign n7820 = n7819 ^ n7569;
  assign n7941 = n7940 ^ n7820;
  assign n7810 = n2102 & n3247;
  assign n7811 = x93 & n2112;
  assign n7812 = x95 & n2381;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = x94 & n2105;
  assign n7815 = n7813 & ~n7814;
  assign n7816 = ~n7810 & n7815;
  assign n7817 = n7816 ^ x26;
  assign n7942 = n7941 ^ n7817;
  assign n7807 = n7689 ^ n7558;
  assign n7808 = ~n7690 & ~n7807;
  assign n7809 = n7808 ^ n7558;
  assign n7943 = n7942 ^ n7809;
  assign n7799 = n1746 & n3763;
  assign n7800 = x96 & n1871;
  assign n7801 = x97 & n1750;
  assign n7802 = ~n7800 & ~n7801;
  assign n7803 = x98 & n1873;
  assign n7804 = n7802 & ~n7803;
  assign n7805 = ~n7799 & n7804;
  assign n7806 = n7805 ^ x23;
  assign n7944 = n7943 ^ n7806;
  assign n7796 = n7691 ^ n7547;
  assign n7797 = n7692 & n7796;
  assign n7798 = n7797 ^ n7547;
  assign n7945 = n7944 ^ n7798;
  assign n7788 = n1404 & n4323;
  assign n7789 = x100 & n1408;
  assign n7790 = x99 & n1514;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = x101 & n1517;
  assign n7793 = n7791 & ~n7792;
  assign n7794 = ~n7788 & n7793;
  assign n7795 = n7794 ^ x20;
  assign n7946 = n7945 ^ n7795;
  assign n7785 = n7693 ^ n7536;
  assign n7786 = ~n7694 & ~n7785;
  assign n7787 = n7786 ^ n7536;
  assign n7947 = n7946 ^ n7787;
  assign n7777 = n1098 & n4912;
  assign n7778 = x103 & n1102;
  assign n7779 = x102 & n1198;
  assign n7780 = ~n7778 & ~n7779;
  assign n7781 = x104 & n1201;
  assign n7782 = n7780 & ~n7781;
  assign n7783 = ~n7777 & n7782;
  assign n7784 = n7783 ^ x17;
  assign n7948 = n7947 ^ n7784;
  assign n7774 = n7695 ^ n7525;
  assign n7775 = n7696 & n7774;
  assign n7776 = n7775 ^ n7525;
  assign n7949 = n7948 ^ n7776;
  assign n7766 = n821 & n5578;
  assign n7767 = x105 & n898;
  assign n7768 = x106 & n824;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = x107 & n901;
  assign n7771 = n7769 & ~n7770;
  assign n7772 = ~n7766 & n7771;
  assign n7773 = n7772 ^ x14;
  assign n7950 = n7949 ^ n7773;
  assign n7763 = n7697 ^ n7506;
  assign n7764 = ~n7698 & ~n7763;
  assign n7765 = n7764 ^ n7506;
  assign n7951 = n7950 ^ n7765;
  assign n7755 = n596 & n6250;
  assign n7756 = x109 & n601;
  assign n7757 = x110 & n676;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = x108 & n673;
  assign n7760 = n7758 & ~n7759;
  assign n7761 = ~n7755 & n7760;
  assign n7762 = n7761 ^ x11;
  assign n7952 = n7951 ^ n7762;
  assign n7750 = n7698 ^ n7506;
  assign n7751 = n7750 ^ n7514;
  assign n7752 = n7514 ^ n7503;
  assign n7753 = n7751 & ~n7752;
  assign n7754 = n7753 ^ n7503;
  assign n7953 = n7952 ^ n7754;
  assign n7742 = n399 & n6975;
  assign n7743 = x111 & n478;
  assign n7744 = x113 & n470;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = x112 & n402;
  assign n7747 = n7745 & ~n7746;
  assign n7748 = ~n7742 & n7747;
  assign n7749 = n7748 ^ x8;
  assign n7954 = n7953 ^ n7749;
  assign n7739 = n7701 ^ n7492;
  assign n7740 = ~n7702 & ~n7739;
  assign n7741 = n7740 ^ n7492;
  assign n7955 = n7954 ^ n7741;
  assign n7730 = n6965 ^ x116;
  assign n7731 = n239 & n7730;
  assign n7732 = x114 & n249;
  assign n7733 = x115 & n242;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = x116 & n280;
  assign n7736 = n7734 & ~n7735;
  assign n7737 = ~n7731 & n7736;
  assign n7738 = n7737 ^ x5;
  assign n7956 = n7955 ^ n7738;
  assign n7727 = n7703 ^ n7480;
  assign n7728 = n7704 & ~n7727;
  assign n7729 = n7728 ^ n7480;
  assign n7957 = n7956 ^ n7729;
  assign n7713 = x118 ^ x117;
  assign n7714 = ~n7464 & n7713;
  assign n7715 = n169 & ~n7714;
  assign n7716 = n7715 ^ x1;
  assign n7717 = n7716 ^ x119;
  assign n7711 = x118 ^ x2;
  assign n7712 = x1 & n7711;
  assign n7718 = n7717 ^ n7712;
  assign n7719 = n7718 ^ n7717;
  assign n7720 = ~x117 & n197;
  assign n7721 = n7720 ^ n7717;
  assign n7722 = n7721 ^ n7717;
  assign n7723 = ~n7719 & ~n7722;
  assign n7724 = n7723 ^ n7717;
  assign n7725 = ~x0 & ~n7724;
  assign n7726 = n7725 ^ n7717;
  assign n7958 = n7957 ^ n7726;
  assign n7708 = n7705 ^ n7460;
  assign n7709 = ~n7706 & n7708;
  assign n7710 = n7709 ^ n7460;
  assign n7959 = n7958 ^ n7710;
  assign n8189 = n420 & n7395;
  assign n8190 = x67 & n7650;
  assign n8191 = x69 & n7652;
  assign n8192 = ~n8190 & ~n8191;
  assign n8193 = x68 & n7400;
  assign n8194 = n8192 & ~n8193;
  assign n8195 = ~n8189 & n8194;
  assign n8196 = n8195 ^ x53;
  assign n8170 = x56 ^ x55;
  assign n8171 = n7644 & n8170;
  assign n8172 = n142 & n8171;
  assign n8173 = x55 & ~n7644;
  assign n8174 = n8173 ^ n7895;
  assign n8175 = ~n8172 & ~n8174;
  assign n8176 = x65 & ~n8175;
  assign n8177 = n7895 ^ x56;
  assign n8178 = n8177 ^ n7895;
  assign n8179 = ~n7644 & n8178;
  assign n8180 = n8179 ^ n7895;
  assign n8181 = n8170 & n8180;
  assign n8182 = x64 & n8181;
  assign n8183 = n152 & n8170;
  assign n8184 = x66 & n7644;
  assign n8185 = ~n8183 & n8184;
  assign n8186 = ~n8182 & ~n8185;
  assign n8187 = ~n8176 & n8186;
  assign n8164 = x55 ^ x53;
  assign n8165 = x64 & n8164;
  assign n8166 = n8165 ^ n233;
  assign n8167 = ~n7644 & ~n8166;
  assign n8168 = n8167 ^ n233;
  assign n8169 = x56 & ~n8168;
  assign n8188 = n8187 ^ n8169;
  assign n8197 = n8196 ^ n8188;
  assign n8161 = n7913 ^ n7910;
  assign n8162 = n7911 & ~n8161;
  assign n8163 = n8162 ^ n7913;
  assign n8198 = n8197 ^ n8163;
  assign n8153 = n575 & n6626;
  assign n8154 = x71 & n6630;
  assign n8155 = x70 & n6884;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = x72 & n6888;
  assign n8158 = n8156 & ~n8157;
  assign n8159 = ~n8153 & n8158;
  assign n8160 = n8159 ^ x50;
  assign n8199 = n8198 ^ n8160;
  assign n8150 = n7914 ^ n7886;
  assign n8151 = ~n7915 & ~n8150;
  assign n8152 = n8151 ^ n7886;
  assign n8200 = n8199 ^ n8152;
  assign n8142 = n789 & n5942;
  assign n8143 = x74 & n5947;
  assign n8144 = x73 & n6186;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = x75 & n6406;
  assign n8147 = n8145 & ~n8146;
  assign n8148 = ~n8142 & n8147;
  assign n8149 = n8148 ^ x47;
  assign n8201 = n8200 ^ n8149;
  assign n8139 = n7916 ^ n7875;
  assign n8140 = n7917 & n8139;
  assign n8141 = n8140 ^ n7875;
  assign n8202 = n8201 ^ n8141;
  assign n8131 = n1041 & n5262;
  assign n8132 = x76 & n5488;
  assign n8133 = x77 & n5266;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = x78 & n5491;
  assign n8136 = n8134 & ~n8135;
  assign n8137 = ~n8131 & n8136;
  assign n8138 = n8137 ^ x44;
  assign n8203 = n8202 ^ n8138;
  assign n8123 = n1340 & n4643;
  assign n8124 = x79 & n4653;
  assign n8125 = x80 & n4646;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = x81 & n5046;
  assign n8128 = n8126 & ~n8127;
  assign n8129 = ~n8123 & n8128;
  assign n8130 = n8129 ^ x41;
  assign n8204 = n8203 ^ n8130;
  assign n8120 = n7929 ^ n7918;
  assign n8121 = ~n7930 & ~n8120;
  assign n8122 = n8121 ^ n7921;
  assign n8205 = n8204 ^ n8122;
  assign n8117 = n7931 ^ n7864;
  assign n8118 = n7932 & n8117;
  assign n8119 = n8118 ^ n7864;
  assign n8206 = n8205 ^ n8119;
  assign n8109 = n1667 & n4040;
  assign n8110 = x82 & n4267;
  assign n8111 = x83 & n4044;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = x84 & n4270;
  assign n8114 = n8112 & ~n8113;
  assign n8115 = ~n8109 & n8114;
  assign n8116 = n8115 ^ x38;
  assign n8207 = n8206 ^ n8116;
  assign n8106 = n7933 ^ n7853;
  assign n8107 = ~n7934 & ~n8106;
  assign n8108 = n8107 ^ n7853;
  assign n8208 = n8207 ^ n8108;
  assign n8098 = n2039 & n3522;
  assign n8099 = x85 & n3699;
  assign n8100 = x86 & n3526;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = x87 & n3701;
  assign n8103 = n8101 & ~n8102;
  assign n8104 = ~n8098 & n8103;
  assign n8105 = n8104 ^ x35;
  assign n8209 = n8208 ^ n8105;
  assign n8095 = n7935 ^ n7842;
  assign n8096 = n7936 & n8095;
  assign n8097 = n8096 ^ n7842;
  assign n8210 = n8209 ^ n8097;
  assign n8087 = n2448 & n3009;
  assign n8088 = x89 & n3013;
  assign n8089 = x88 & n3181;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = x90 & n3183;
  assign n8092 = n8090 & ~n8091;
  assign n8093 = ~n8087 & n8092;
  assign n8094 = n8093 ^ x32;
  assign n8211 = n8210 ^ n8094;
  assign n8084 = n7937 ^ n7831;
  assign n8085 = ~n7938 & ~n8084;
  assign n8086 = n8085 ^ n7831;
  assign n8212 = n8211 ^ n8086;
  assign n8076 = n2527 & n2901;
  assign n8077 = x91 & n2690;
  assign n8078 = x92 & n2530;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = x93 & n2693;
  assign n8081 = n8079 & ~n8080;
  assign n8082 = ~n8076 & n8081;
  assign n8083 = n8082 ^ x29;
  assign n8213 = n8212 ^ n8083;
  assign n8073 = n7939 ^ n7820;
  assign n8074 = n7940 & n8073;
  assign n8075 = n8074 ^ n7820;
  assign n8214 = n8213 ^ n8075;
  assign n8065 = n2102 & n3403;
  assign n8066 = x94 & n2112;
  assign n8067 = x95 & n2105;
  assign n8068 = ~n8066 & ~n8067;
  assign n8069 = x96 & n2381;
  assign n8070 = n8068 & ~n8069;
  assign n8071 = ~n8065 & n8070;
  assign n8072 = n8071 ^ x26;
  assign n8215 = n8214 ^ n8072;
  assign n8062 = n7941 ^ n7809;
  assign n8063 = ~n7942 & ~n8062;
  assign n8064 = n8063 ^ n7809;
  assign n8216 = n8215 ^ n8064;
  assign n8054 = n1746 & n3943;
  assign n8055 = x97 & n1871;
  assign n8056 = x98 & n1750;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = x99 & n1873;
  assign n8059 = n8057 & ~n8058;
  assign n8060 = ~n8054 & n8059;
  assign n8061 = n8060 ^ x23;
  assign n8217 = n8216 ^ n8061;
  assign n8051 = n7943 ^ n7798;
  assign n8052 = n7944 & n8051;
  assign n8053 = n8052 ^ n7798;
  assign n8218 = n8217 ^ n8053;
  assign n8043 = n1404 & n4509;
  assign n8044 = x100 & n1514;
  assign n8045 = x101 & n1408;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = x102 & n1517;
  assign n8048 = n8046 & ~n8047;
  assign n8049 = ~n8043 & n8048;
  assign n8050 = n8049 ^ x20;
  assign n8219 = n8218 ^ n8050;
  assign n8040 = n7945 ^ n7787;
  assign n8041 = ~n7946 & ~n8040;
  assign n8042 = n8041 ^ n7787;
  assign n8220 = n8219 ^ n8042;
  assign n8032 = n1098 & n5117;
  assign n8033 = x103 & n1198;
  assign n8034 = x104 & n1102;
  assign n8035 = ~n8033 & ~n8034;
  assign n8036 = x105 & n1201;
  assign n8037 = n8035 & ~n8036;
  assign n8038 = ~n8032 & n8037;
  assign n8039 = n8038 ^ x17;
  assign n8221 = n8220 ^ n8039;
  assign n8029 = n7947 ^ n7776;
  assign n8030 = n7948 & n8029;
  assign n8031 = n8030 ^ n7776;
  assign n8222 = n8221 ^ n8031;
  assign n8021 = n821 & n5792;
  assign n8022 = x106 & n898;
  assign n8023 = x107 & n824;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = x108 & n901;
  assign n8026 = n8024 & ~n8025;
  assign n8027 = ~n8021 & n8026;
  assign n8028 = n8027 ^ x14;
  assign n8223 = n8222 ^ n8028;
  assign n8018 = n7949 ^ n7765;
  assign n8019 = ~n7950 & ~n8018;
  assign n8020 = n8019 ^ n7765;
  assign n8224 = n8223 ^ n8020;
  assign n8010 = n596 & n6478;
  assign n8011 = x109 & n673;
  assign n8012 = x111 & n676;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = x110 & n601;
  assign n8015 = n8013 & ~n8014;
  assign n8016 = ~n8010 & n8015;
  assign n8017 = n8016 ^ x11;
  assign n8225 = n8224 ^ n8017;
  assign n8007 = n7951 ^ n7754;
  assign n8008 = n7952 & n8007;
  assign n8009 = n8008 ^ n7754;
  assign n8226 = n8225 ^ n8009;
  assign n7999 = n399 & n7220;
  assign n8000 = x112 & n478;
  assign n8001 = x113 & n402;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = x114 & n470;
  assign n8004 = n8002 & ~n8003;
  assign n8005 = ~n7999 & n8004;
  assign n8006 = n8005 ^ x8;
  assign n8227 = n8226 ^ n8006;
  assign n7996 = n7953 ^ n7741;
  assign n7997 = ~n7954 & ~n7996;
  assign n7998 = n7997 ^ n7741;
  assign n8228 = n8227 ^ n7998;
  assign n7987 = n7210 ^ x117;
  assign n7988 = n239 & n7987;
  assign n7989 = x115 & n249;
  assign n7990 = x116 & n242;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = x117 & n280;
  assign n7993 = n7991 & ~n7992;
  assign n7994 = ~n7988 & n7993;
  assign n7995 = n7994 ^ x5;
  assign n8229 = n8228 ^ n7995;
  assign n7984 = n7955 ^ n7729;
  assign n7985 = n7956 & ~n7984;
  assign n7986 = n7985 ^ n7729;
  assign n8230 = n8229 ^ n7986;
  assign n7964 = x119 ^ x118;
  assign n7965 = n7463 ^ n7462;
  assign n7966 = n7462 ^ x119;
  assign n7967 = n7966 ^ n7462;
  assign n7968 = n7965 & ~n7967;
  assign n7969 = n7968 ^ n7462;
  assign n7970 = n7964 & ~n7969;
  assign n7971 = n169 & ~n7970;
  assign n7972 = n7971 ^ x1;
  assign n7973 = n7972 ^ x120;
  assign n7963 = ~x118 & n197;
  assign n7974 = n7973 ^ n7963;
  assign n7975 = n7974 ^ n7973;
  assign n7976 = x119 ^ x2;
  assign n7977 = x1 & n7976;
  assign n7978 = n7977 ^ n7973;
  assign n7979 = n7978 ^ n7973;
  assign n7980 = ~n7975 & ~n7979;
  assign n7981 = n7980 ^ n7973;
  assign n7982 = ~x0 & ~n7981;
  assign n7983 = n7982 ^ n7973;
  assign n8231 = n8230 ^ n7983;
  assign n7960 = n7957 ^ n7710;
  assign n7961 = ~n7958 & n7960;
  assign n7962 = n7961 ^ n7710;
  assign n8232 = n8231 ^ n7962;
  assign n8479 = n1149 & n5262;
  assign n8480 = x77 & n5488;
  assign n8481 = x79 & n5491;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = x78 & n5266;
  assign n8484 = n8482 & ~n8483;
  assign n8485 = ~n8479 & n8484;
  assign n8486 = n8485 ^ x44;
  assign n8476 = n8202 ^ n8122;
  assign n8477 = n8203 & n8476;
  assign n8478 = n8477 ^ n8122;
  assign n8487 = n8486 ^ n8478;
  assign n8464 = ~n653 & n6626;
  assign n8465 = x72 & n6630;
  assign n8466 = x71 & n6884;
  assign n8467 = ~n8465 & ~n8466;
  assign n8468 = x73 & n6888;
  assign n8469 = n8467 & ~n8468;
  assign n8470 = ~n8464 & n8469;
  assign n8471 = n8470 ^ x50;
  assign n8461 = n8198 ^ n8152;
  assign n8462 = n8199 & n8461;
  assign n8463 = n8462 ^ n8152;
  assign n8472 = n8471 ^ n8463;
  assign n8451 = n458 & n7395;
  assign n8452 = x68 & n7650;
  assign n8453 = x69 & n7400;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = x70 & n7652;
  assign n8456 = n8454 & ~n8455;
  assign n8457 = ~n8451 & n8456;
  assign n8458 = n8457 ^ x53;
  assign n8448 = n8196 ^ n8163;
  assign n8449 = ~n8197 & ~n8448;
  assign n8450 = n8449 ^ n8163;
  assign n8459 = n8458 ^ n8450;
  assign n8417 = n168 & n8170;
  assign n8418 = n8417 ^ x67;
  assign n8419 = n7644 & n8418;
  assign n8420 = x65 & n8181;
  assign n8421 = x66 & n8174;
  assign n8422 = ~n8420 & ~n8421;
  assign n8423 = ~n8419 & n8422;
  assign n8424 = n8423 ^ x56;
  assign n8425 = x56 & n8168;
  assign n8436 = n8187 & n8425;
  assign n8427 = x57 ^ x56;
  assign n8437 = x64 & n8427;
  assign n8438 = ~n8436 & ~n8437;
  assign n8426 = n8187 ^ x57;
  assign n8428 = n8427 ^ n8426;
  assign n8429 = n8428 ^ n8427;
  assign n8430 = n8427 ^ x64;
  assign n8431 = n8430 ^ n8427;
  assign n8432 = n8429 & n8431;
  assign n8433 = n8432 ^ n8427;
  assign n8434 = n8425 & ~n8433;
  assign n8435 = n8434 ^ n8427;
  assign n8439 = n8438 ^ n8435;
  assign n8440 = n8439 ^ n8438;
  assign n8441 = ~x64 & ~n8436;
  assign n8442 = n8441 ^ n8438;
  assign n8443 = n8442 ^ n8438;
  assign n8444 = n8440 & ~n8443;
  assign n8445 = n8444 ^ n8438;
  assign n8446 = ~n8424 & n8445;
  assign n8447 = n8446 ^ n8438;
  assign n8460 = n8459 ^ n8447;
  assign n8473 = n8472 ^ n8460;
  assign n8409 = n870 & n5942;
  assign n8410 = x74 & n6186;
  assign n8411 = x76 & n6406;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = x75 & n5947;
  assign n8414 = n8412 & ~n8413;
  assign n8415 = ~n8409 & n8414;
  assign n8416 = n8415 ^ x47;
  assign n8474 = n8473 ^ n8416;
  assign n8406 = n8200 ^ n8141;
  assign n8407 = ~n8201 & ~n8406;
  assign n8408 = n8407 ^ n8141;
  assign n8475 = n8474 ^ n8408;
  assign n8488 = n8487 ^ n8475;
  assign n8398 = n1454 & n4643;
  assign n8399 = x80 & n4653;
  assign n8400 = x81 & n4646;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = x82 & n5046;
  assign n8403 = n8401 & ~n8402;
  assign n8404 = ~n8398 & n8403;
  assign n8405 = n8404 ^ x41;
  assign n8489 = n8488 ^ n8405;
  assign n8395 = n8130 ^ n8119;
  assign n8396 = ~n8205 & ~n8395;
  assign n8397 = n8396 ^ n8119;
  assign n8490 = n8489 ^ n8397;
  assign n8387 = n1801 & n4040;
  assign n8388 = x83 & n4267;
  assign n8389 = x85 & n4270;
  assign n8390 = ~n8388 & ~n8389;
  assign n8391 = x84 & n4044;
  assign n8392 = n8390 & ~n8391;
  assign n8393 = ~n8387 & n8392;
  assign n8394 = n8393 ^ x38;
  assign n8491 = n8490 ^ n8394;
  assign n8384 = n8206 ^ n8108;
  assign n8385 = n8207 & n8384;
  assign n8386 = n8385 ^ n8108;
  assign n8492 = n8491 ^ n8386;
  assign n8376 = n2176 & n3522;
  assign n8377 = x86 & n3699;
  assign n8378 = x87 & n3526;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = x88 & n3701;
  assign n8381 = n8379 & ~n8380;
  assign n8382 = ~n8376 & n8381;
  assign n8383 = n8382 ^ x35;
  assign n8493 = n8492 ^ n8383;
  assign n8373 = n8208 ^ n8097;
  assign n8374 = ~n8209 & ~n8373;
  assign n8375 = n8374 ^ n8097;
  assign n8494 = n8493 ^ n8375;
  assign n8365 = n2607 & n3009;
  assign n8366 = x89 & n3181;
  assign n8367 = x90 & n3013;
  assign n8368 = ~n8366 & ~n8367;
  assign n8369 = x91 & n3183;
  assign n8370 = n8368 & ~n8369;
  assign n8371 = ~n8365 & n8370;
  assign n8372 = n8371 ^ x32;
  assign n8495 = n8494 ^ n8372;
  assign n8362 = n8210 ^ n8086;
  assign n8363 = n8211 & n8362;
  assign n8364 = n8363 ^ n8086;
  assign n8496 = n8495 ^ n8364;
  assign n8354 = n2527 & n3078;
  assign n8355 = x92 & n2690;
  assign n8356 = x93 & n2530;
  assign n8357 = ~n8355 & ~n8356;
  assign n8358 = x94 & n2693;
  assign n8359 = n8357 & ~n8358;
  assign n8360 = ~n8354 & n8359;
  assign n8361 = n8360 ^ x29;
  assign n8497 = n8496 ^ n8361;
  assign n8351 = n8212 ^ n8075;
  assign n8352 = ~n8213 & ~n8351;
  assign n8353 = n8352 ^ n8075;
  assign n8498 = n8497 ^ n8353;
  assign n8343 = n2102 & n3585;
  assign n8344 = x95 & n2112;
  assign n8345 = x97 & n2381;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = x96 & n2105;
  assign n8348 = n8346 & ~n8347;
  assign n8349 = ~n8343 & n8348;
  assign n8350 = n8349 ^ x26;
  assign n8499 = n8498 ^ n8350;
  assign n8340 = n8214 ^ n8064;
  assign n8341 = n8215 & n8340;
  assign n8342 = n8341 ^ n8064;
  assign n8500 = n8499 ^ n8342;
  assign n8332 = n1746 & n4141;
  assign n8333 = x98 & n1871;
  assign n8334 = x99 & n1750;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = x100 & n1873;
  assign n8337 = n8335 & ~n8336;
  assign n8338 = ~n8332 & n8337;
  assign n8339 = n8338 ^ x23;
  assign n8501 = n8500 ^ n8339;
  assign n8329 = n8216 ^ n8053;
  assign n8330 = ~n8217 & ~n8329;
  assign n8331 = n8330 ^ n8053;
  assign n8502 = n8501 ^ n8331;
  assign n8321 = n1404 & n4718;
  assign n8322 = x101 & n1514;
  assign n8323 = x103 & n1517;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = x102 & n1408;
  assign n8326 = n8324 & ~n8325;
  assign n8327 = ~n8321 & n8326;
  assign n8328 = n8327 ^ x20;
  assign n8503 = n8502 ^ n8328;
  assign n8318 = n8218 ^ n8042;
  assign n8319 = n8219 & n8318;
  assign n8320 = n8319 ^ n8042;
  assign n8504 = n8503 ^ n8320;
  assign n8310 = n1098 & n5351;
  assign n8311 = x104 & n1198;
  assign n8312 = x105 & n1102;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = x106 & n1201;
  assign n8315 = n8313 & ~n8314;
  assign n8316 = ~n8310 & n8315;
  assign n8317 = n8316 ^ x17;
  assign n8505 = n8504 ^ n8317;
  assign n8307 = n8220 ^ n8031;
  assign n8308 = ~n8221 & ~n8307;
  assign n8309 = n8308 ^ n8031;
  assign n8506 = n8505 ^ n8309;
  assign n8299 = n821 & n6026;
  assign n8300 = x107 & n898;
  assign n8301 = x108 & n824;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = x109 & n901;
  assign n8304 = n8302 & ~n8303;
  assign n8305 = ~n8299 & n8304;
  assign n8306 = n8305 ^ x14;
  assign n8507 = n8506 ^ n8306;
  assign n8296 = n8222 ^ n8020;
  assign n8297 = n8223 & n8296;
  assign n8298 = n8297 ^ n8020;
  assign n8508 = n8507 ^ n8298;
  assign n8288 = n596 & n6728;
  assign n8289 = x110 & n673;
  assign n8290 = x112 & n676;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = x111 & n601;
  assign n8293 = n8291 & ~n8292;
  assign n8294 = ~n8288 & n8293;
  assign n8295 = n8294 ^ x11;
  assign n8509 = n8508 ^ n8295;
  assign n8285 = n8224 ^ n8009;
  assign n8286 = ~n8225 & ~n8285;
  assign n8287 = n8286 ^ n8009;
  assign n8510 = n8509 ^ n8287;
  assign n8277 = n399 & n7481;
  assign n8278 = x113 & n478;
  assign n8279 = x114 & n402;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = x115 & n470;
  assign n8282 = n8280 & ~n8281;
  assign n8283 = ~n8277 & n8282;
  assign n8284 = n8283 ^ x8;
  assign n8511 = n8510 ^ n8284;
  assign n8274 = n8226 ^ n7998;
  assign n8275 = n8227 & n8274;
  assign n8276 = n8275 ^ n7998;
  assign n8512 = n8511 ^ n8276;
  assign n8238 = ~n7208 & ~n7463;
  assign n8265 = n8238 ^ n7713;
  assign n8266 = n239 & n8265;
  assign n8267 = x116 & n249;
  assign n8268 = x118 & n280;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = x117 & n242;
  assign n8271 = n8269 & ~n8270;
  assign n8272 = ~n8266 & n8271;
  assign n8273 = n8272 ^ x5;
  assign n8513 = n8512 ^ n8273;
  assign n8262 = n8228 ^ n7986;
  assign n8263 = ~n8229 & n8262;
  assign n8264 = n8263 ^ n7986;
  assign n8514 = n8513 ^ n8264;
  assign n8239 = ~x118 & ~x120;
  assign n8240 = ~x117 & ~x119;
  assign n8241 = ~n8239 & ~n8240;
  assign n8242 = ~n8238 & ~n8241;
  assign n8243 = ~x117 & n8239;
  assign n8244 = ~x119 & x120;
  assign n8245 = x118 & n8244;
  assign n8246 = n8245 ^ x119;
  assign n8247 = ~n8243 & n8246;
  assign n8248 = ~n8242 & n8247;
  assign n8249 = n8248 ^ x120;
  assign n8250 = n169 & ~n8249;
  assign n8251 = n8250 ^ x1;
  assign n8252 = n8251 ^ x121;
  assign n8236 = x120 ^ x2;
  assign n8237 = x1 & n8236;
  assign n8253 = n8252 ^ n8237;
  assign n8254 = n8253 ^ n8252;
  assign n8255 = ~x119 & n197;
  assign n8256 = n8255 ^ n8252;
  assign n8257 = n8256 ^ n8252;
  assign n8258 = ~n8254 & ~n8257;
  assign n8259 = n8258 ^ n8252;
  assign n8260 = ~x0 & ~n8259;
  assign n8261 = n8260 ^ n8252;
  assign n8515 = n8514 ^ n8261;
  assign n8233 = n8230 ^ n7962;
  assign n8234 = n8231 & ~n8233;
  assign n8235 = n8234 ^ n7962;
  assign n8516 = n8515 ^ n8235;
  assign n8742 = x56 & x57;
  assign n8743 = n8742 ^ x58;
  assign n8744 = ~x64 & n8743;
  assign n8738 = x65 ^ x57;
  assign n8739 = n8427 & ~n8738;
  assign n8740 = n8739 ^ x56;
  assign n8741 = n8740 ^ x58;
  assign n8745 = n8744 ^ n8741;
  assign n8737 = ~n8424 & ~n8438;
  assign n8746 = n8745 ^ n8737;
  assign n8728 = n321 & n8171;
  assign n8729 = x67 & n8174;
  assign n8730 = x66 & n8181;
  assign n8731 = ~n8729 & ~n8730;
  assign n8732 = n7644 & ~n8170;
  assign n8733 = x68 & n8732;
  assign n8734 = n8731 & ~n8733;
  assign n8735 = ~n8728 & n8734;
  assign n8736 = n8735 ^ x56;
  assign n8747 = n8746 ^ n8736;
  assign n8720 = n517 & n7395;
  assign n8721 = x70 & n7400;
  assign n8722 = x69 & n7650;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = x71 & n7652;
  assign n8725 = n8723 & ~n8724;
  assign n8726 = ~n8720 & n8725;
  assign n8727 = n8726 ^ x53;
  assign n8748 = n8747 ^ n8727;
  assign n8717 = n8458 ^ n8447;
  assign n8718 = ~n8459 & ~n8717;
  assign n8719 = n8718 ^ n8450;
  assign n8749 = n8748 ^ n8719;
  assign n8709 = ~n721 & n6626;
  assign n8710 = x73 & n6630;
  assign n8711 = x72 & n6884;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = x74 & n6888;
  assign n8714 = n8712 & ~n8713;
  assign n8715 = ~n8709 & n8714;
  assign n8716 = n8715 ^ x50;
  assign n8750 = n8749 ^ n8716;
  assign n8706 = n8471 ^ n8460;
  assign n8707 = ~n8472 & n8706;
  assign n8708 = n8707 ^ n8463;
  assign n8751 = n8750 ^ n8708;
  assign n8698 = n956 & n5942;
  assign n8699 = x75 & n6186;
  assign n8700 = x76 & n5947;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = x77 & n6406;
  assign n8703 = n8701 & ~n8702;
  assign n8704 = ~n8698 & n8703;
  assign n8705 = n8704 ^ x47;
  assign n8752 = n8751 ^ n8705;
  assign n8695 = n8473 ^ n8408;
  assign n8696 = ~n8474 & ~n8695;
  assign n8697 = n8696 ^ n8408;
  assign n8753 = n8752 ^ n8697;
  assign n8687 = n1242 & n5262;
  assign n8688 = x79 & n5266;
  assign n8689 = x80 & n5491;
  assign n8690 = ~n8688 & ~n8689;
  assign n8691 = x78 & n5488;
  assign n8692 = n8690 & ~n8691;
  assign n8693 = ~n8687 & n8692;
  assign n8694 = n8693 ^ x44;
  assign n8754 = n8753 ^ n8694;
  assign n8684 = n8486 ^ n8475;
  assign n8685 = ~n8487 & n8684;
  assign n8686 = n8685 ^ n8478;
  assign n8755 = n8754 ^ n8686;
  assign n8676 = n1560 & n4643;
  assign n8677 = x81 & n4653;
  assign n8678 = x82 & n4646;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = x83 & n5046;
  assign n8681 = n8679 & ~n8680;
  assign n8682 = ~n8676 & n8681;
  assign n8683 = n8682 ^ x41;
  assign n8756 = n8755 ^ n8683;
  assign n8673 = n8488 ^ n8397;
  assign n8674 = ~n8489 & ~n8673;
  assign n8675 = n8674 ^ n8397;
  assign n8757 = n8756 ^ n8675;
  assign n8665 = n1920 & n4040;
  assign n8666 = x84 & n4267;
  assign n8667 = x86 & n4270;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = x85 & n4044;
  assign n8670 = n8668 & ~n8669;
  assign n8671 = ~n8665 & n8670;
  assign n8672 = n8671 ^ x38;
  assign n8758 = n8757 ^ n8672;
  assign n8662 = n8490 ^ n8386;
  assign n8663 = n8491 & n8662;
  assign n8664 = n8663 ^ n8386;
  assign n8759 = n8758 ^ n8664;
  assign n8654 = n2310 & n3522;
  assign n8655 = x87 & n3699;
  assign n8656 = x89 & n3701;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = x88 & n3526;
  assign n8659 = n8657 & ~n8658;
  assign n8660 = ~n8654 & n8659;
  assign n8661 = n8660 ^ x35;
  assign n8760 = n8759 ^ n8661;
  assign n8651 = n8492 ^ n8375;
  assign n8652 = ~n8493 & ~n8651;
  assign n8653 = n8652 ^ n8375;
  assign n8761 = n8760 ^ n8653;
  assign n8643 = n2755 & n3009;
  assign n8644 = x91 & n3013;
  assign n8645 = x90 & n3181;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = x92 & n3183;
  assign n8648 = n8646 & ~n8647;
  assign n8649 = ~n8643 & n8648;
  assign n8650 = n8649 ^ x32;
  assign n8762 = n8761 ^ n8650;
  assign n8640 = n8494 ^ n8364;
  assign n8641 = n8495 & n8640;
  assign n8642 = n8641 ^ n8364;
  assign n8763 = n8762 ^ n8642;
  assign n8632 = n2527 & n3247;
  assign n8633 = x93 & n2690;
  assign n8634 = x94 & n2530;
  assign n8635 = ~n8633 & ~n8634;
  assign n8636 = x95 & n2693;
  assign n8637 = n8635 & ~n8636;
  assign n8638 = ~n8632 & n8637;
  assign n8639 = n8638 ^ x29;
  assign n8764 = n8763 ^ n8639;
  assign n8629 = n8496 ^ n8353;
  assign n8630 = ~n8497 & ~n8629;
  assign n8631 = n8630 ^ n8353;
  assign n8765 = n8764 ^ n8631;
  assign n8621 = n2102 & n3763;
  assign n8622 = x96 & n2112;
  assign n8623 = x97 & n2105;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = x98 & n2381;
  assign n8626 = n8624 & ~n8625;
  assign n8627 = ~n8621 & n8626;
  assign n8628 = n8627 ^ x26;
  assign n8766 = n8765 ^ n8628;
  assign n8618 = n8498 ^ n8342;
  assign n8619 = n8499 & n8618;
  assign n8620 = n8619 ^ n8342;
  assign n8767 = n8766 ^ n8620;
  assign n8610 = n1746 & n4323;
  assign n8611 = x100 & n1750;
  assign n8612 = x99 & n1871;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = x101 & n1873;
  assign n8615 = n8613 & ~n8614;
  assign n8616 = ~n8610 & n8615;
  assign n8617 = n8616 ^ x23;
  assign n8768 = n8767 ^ n8617;
  assign n8607 = n8500 ^ n8331;
  assign n8608 = ~n8501 & ~n8607;
  assign n8609 = n8608 ^ n8331;
  assign n8769 = n8768 ^ n8609;
  assign n8599 = n1404 & n4912;
  assign n8600 = x102 & n1514;
  assign n8601 = x103 & n1408;
  assign n8602 = ~n8600 & ~n8601;
  assign n8603 = x104 & n1517;
  assign n8604 = n8602 & ~n8603;
  assign n8605 = ~n8599 & n8604;
  assign n8606 = n8605 ^ x20;
  assign n8770 = n8769 ^ n8606;
  assign n8596 = n8502 ^ n8320;
  assign n8597 = n8503 & n8596;
  assign n8598 = n8597 ^ n8320;
  assign n8771 = n8770 ^ n8598;
  assign n8588 = n1098 & n5578;
  assign n8589 = x105 & n1198;
  assign n8590 = x106 & n1102;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = x107 & n1201;
  assign n8593 = n8591 & ~n8592;
  assign n8594 = ~n8588 & n8593;
  assign n8595 = n8594 ^ x17;
  assign n8772 = n8771 ^ n8595;
  assign n8585 = n8504 ^ n8309;
  assign n8586 = ~n8505 & ~n8585;
  assign n8587 = n8586 ^ n8309;
  assign n8773 = n8772 ^ n8587;
  assign n8577 = n821 & n6250;
  assign n8578 = x108 & n898;
  assign n8579 = x109 & n824;
  assign n8580 = ~n8578 & ~n8579;
  assign n8581 = x110 & n901;
  assign n8582 = n8580 & ~n8581;
  assign n8583 = ~n8577 & n8582;
  assign n8584 = n8583 ^ x14;
  assign n8774 = n8773 ^ n8584;
  assign n8574 = n8506 ^ n8298;
  assign n8575 = n8507 & n8574;
  assign n8576 = n8575 ^ n8298;
  assign n8775 = n8774 ^ n8576;
  assign n8566 = n596 & n6975;
  assign n8567 = x111 & n673;
  assign n8568 = x112 & n601;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = x113 & n676;
  assign n8571 = n8569 & ~n8570;
  assign n8572 = ~n8566 & n8571;
  assign n8573 = n8572 ^ x11;
  assign n8776 = n8775 ^ n8573;
  assign n8563 = n8508 ^ n8287;
  assign n8564 = ~n8509 & ~n8563;
  assign n8565 = n8564 ^ n8287;
  assign n8777 = n8776 ^ n8565;
  assign n8555 = n399 & n7730;
  assign n8556 = x114 & n478;
  assign n8557 = x115 & n402;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = x116 & n470;
  assign n8560 = n8558 & ~n8559;
  assign n8561 = ~n8555 & n8560;
  assign n8562 = n8561 ^ x8;
  assign n8778 = n8777 ^ n8562;
  assign n8552 = n8510 ^ n8276;
  assign n8553 = n8511 & n8552;
  assign n8554 = n8553 ^ n8276;
  assign n8779 = n8778 ^ n8554;
  assign n8542 = n7714 ^ x119;
  assign n8543 = n239 & n8542;
  assign n8544 = x117 & n249;
  assign n8545 = x119 & n280;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = x118 & n242;
  assign n8548 = n8546 & ~n8547;
  assign n8549 = ~n8543 & n8548;
  assign n8550 = n8549 ^ x5;
  assign n8524 = x120 & n8248;
  assign n8525 = ~x121 & ~n8524;
  assign n8526 = ~x120 & ~n8248;
  assign n8527 = x121 & ~n8526;
  assign n8528 = ~n8525 & ~n8527;
  assign n8529 = n169 & ~n8528;
  assign n8530 = n8529 ^ x1;
  assign n8531 = n8530 ^ x122;
  assign n8523 = ~x120 & n197;
  assign n8532 = n8531 ^ n8523;
  assign n8533 = n8532 ^ n8531;
  assign n8534 = x121 ^ x2;
  assign n8535 = x1 & n8534;
  assign n8536 = n8535 ^ n8531;
  assign n8537 = n8536 ^ n8531;
  assign n8538 = ~n8533 & ~n8537;
  assign n8539 = n8538 ^ n8531;
  assign n8540 = ~x0 & ~n8539;
  assign n8541 = n8540 ^ n8531;
  assign n8551 = n8550 ^ n8541;
  assign n8780 = n8779 ^ n8551;
  assign n8520 = n8512 ^ n8264;
  assign n8521 = ~n8513 & n8520;
  assign n8522 = n8521 ^ n8264;
  assign n8781 = n8780 ^ n8522;
  assign n8517 = n8514 ^ n8235;
  assign n8518 = n8515 & ~n8517;
  assign n8519 = n8518 ^ n8235;
  assign n8782 = n8781 ^ n8519;
  assign n9040 = n1041 & n5942;
  assign n9041 = x77 & n5947;
  assign n9042 = x76 & n6186;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = x78 & n6406;
  assign n9045 = n9043 & ~n9044;
  assign n9046 = ~n9040 & n9045;
  assign n9047 = n9046 ^ x47;
  assign n9037 = n8751 ^ n8697;
  assign n9038 = ~n8752 & ~n9037;
  assign n9039 = n9038 ^ n8697;
  assign n9048 = n9047 ^ n9039;
  assign n9027 = n789 & n6626;
  assign n9028 = x73 & n6884;
  assign n9029 = x75 & n6888;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = x74 & n6630;
  assign n9032 = n9030 & ~n9031;
  assign n9033 = ~n9027 & n9032;
  assign n9034 = n9033 ^ x50;
  assign n9024 = n8749 ^ n8708;
  assign n9025 = n8750 & n9024;
  assign n9026 = n9025 ^ n8708;
  assign n9035 = n9034 ^ n9026;
  assign n9001 = x59 ^ x58;
  assign n9002 = n8427 & n9001;
  assign n9003 = n142 & n9002;
  assign n9004 = x58 & ~n8427;
  assign n9005 = n9004 ^ n8742;
  assign n9006 = ~n9003 & ~n9005;
  assign n9007 = x65 & ~n9006;
  assign n9008 = n8742 ^ x59;
  assign n9009 = n9008 ^ n8742;
  assign n9010 = ~n8427 & n9009;
  assign n9011 = n9010 ^ n8742;
  assign n9012 = n9001 & n9011;
  assign n9013 = x64 & n9012;
  assign n9014 = n152 & n9001;
  assign n9015 = x66 & n8427;
  assign n9016 = ~n9014 & n9015;
  assign n9017 = ~n9013 & ~n9016;
  assign n9018 = ~n9007 & n9017;
  assign n8995 = x58 ^ x56;
  assign n8996 = x64 & n8995;
  assign n8997 = n8996 ^ n233;
  assign n8998 = ~n8427 & ~n8997;
  assign n8999 = n8998 ^ n233;
  assign n9000 = x59 & ~n8999;
  assign n9019 = n9018 ^ n9000;
  assign n8992 = n8745 ^ n8736;
  assign n8993 = n8746 & n8992;
  assign n8994 = n8993 ^ n8737;
  assign n9020 = n9019 ^ n8994;
  assign n8984 = n420 & n8171;
  assign n8985 = x68 & n8174;
  assign n8986 = x67 & n8181;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = x69 & n8732;
  assign n8989 = n8987 & ~n8988;
  assign n8990 = ~n8984 & n8989;
  assign n8991 = n8990 ^ x56;
  assign n9021 = n9020 ^ n8991;
  assign n8976 = n575 & n7395;
  assign n8977 = x70 & n7650;
  assign n8978 = x72 & n7652;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = x71 & n7400;
  assign n8981 = n8979 & ~n8980;
  assign n8982 = ~n8976 & n8981;
  assign n8983 = n8982 ^ x53;
  assign n9022 = n9021 ^ n8983;
  assign n8973 = n8747 ^ n8719;
  assign n8974 = ~n8748 & ~n8973;
  assign n8975 = n8974 ^ n8719;
  assign n9023 = n9022 ^ n8975;
  assign n9036 = n9035 ^ n9023;
  assign n9049 = n9048 ^ n9036;
  assign n8965 = n1340 & n5262;
  assign n8966 = x79 & n5488;
  assign n8967 = x80 & n5266;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = x81 & n5491;
  assign n8970 = n8968 & ~n8969;
  assign n8971 = ~n8965 & n8970;
  assign n8972 = n8971 ^ x44;
  assign n9050 = n9049 ^ n8972;
  assign n8962 = n8753 ^ n8686;
  assign n8963 = n8754 & n8962;
  assign n8964 = n8963 ^ n8686;
  assign n9051 = n9050 ^ n8964;
  assign n8954 = n1667 & n4643;
  assign n8955 = x82 & n4653;
  assign n8956 = x83 & n4646;
  assign n8957 = ~n8955 & ~n8956;
  assign n8958 = x84 & n5046;
  assign n8959 = n8957 & ~n8958;
  assign n8960 = ~n8954 & n8959;
  assign n8961 = n8960 ^ x41;
  assign n9052 = n9051 ^ n8961;
  assign n8951 = n8755 ^ n8675;
  assign n8952 = ~n8756 & ~n8951;
  assign n8953 = n8952 ^ n8675;
  assign n9053 = n9052 ^ n8953;
  assign n8943 = n2039 & n4040;
  assign n8944 = x85 & n4267;
  assign n8945 = x86 & n4044;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = x87 & n4270;
  assign n8948 = n8946 & ~n8947;
  assign n8949 = ~n8943 & n8948;
  assign n8950 = n8949 ^ x38;
  assign n9054 = n9053 ^ n8950;
  assign n8940 = n8757 ^ n8664;
  assign n8941 = n8758 & n8940;
  assign n8942 = n8941 ^ n8664;
  assign n9055 = n9054 ^ n8942;
  assign n8932 = n2448 & n3522;
  assign n8933 = x88 & n3699;
  assign n8934 = x90 & n3701;
  assign n8935 = ~n8933 & ~n8934;
  assign n8936 = x89 & n3526;
  assign n8937 = n8935 & ~n8936;
  assign n8938 = ~n8932 & n8937;
  assign n8939 = n8938 ^ x35;
  assign n9056 = n9055 ^ n8939;
  assign n8929 = n8759 ^ n8653;
  assign n8930 = ~n8760 & ~n8929;
  assign n8931 = n8930 ^ n8653;
  assign n9057 = n9056 ^ n8931;
  assign n8921 = n2901 & n3009;
  assign n8922 = x92 & n3013;
  assign n8923 = x91 & n3181;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = x93 & n3183;
  assign n8926 = n8924 & ~n8925;
  assign n8927 = ~n8921 & n8926;
  assign n8928 = n8927 ^ x32;
  assign n9058 = n9057 ^ n8928;
  assign n8918 = n8761 ^ n8642;
  assign n8919 = n8762 & n8918;
  assign n8920 = n8919 ^ n8642;
  assign n9059 = n9058 ^ n8920;
  assign n8910 = n2527 & n3403;
  assign n8911 = x94 & n2690;
  assign n8912 = x95 & n2530;
  assign n8913 = ~n8911 & ~n8912;
  assign n8914 = x96 & n2693;
  assign n8915 = n8913 & ~n8914;
  assign n8916 = ~n8910 & n8915;
  assign n8917 = n8916 ^ x29;
  assign n9060 = n9059 ^ n8917;
  assign n8907 = n8639 ^ n8631;
  assign n8908 = n8764 & n8907;
  assign n8909 = n8908 ^ n8763;
  assign n9061 = n9060 ^ n8909;
  assign n8899 = n2102 & n3943;
  assign n8900 = x97 & n2112;
  assign n8901 = x99 & n2381;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = x98 & n2105;
  assign n8904 = n8902 & ~n8903;
  assign n8905 = ~n8899 & n8904;
  assign n8906 = n8905 ^ x26;
  assign n9062 = n9061 ^ n8906;
  assign n8896 = n8765 ^ n8620;
  assign n8897 = n8766 & n8896;
  assign n8898 = n8897 ^ n8620;
  assign n9063 = n9062 ^ n8898;
  assign n8888 = n1746 & n4509;
  assign n8889 = x100 & n1871;
  assign n8890 = x101 & n1750;
  assign n8891 = ~n8889 & ~n8890;
  assign n8892 = x102 & n1873;
  assign n8893 = n8891 & ~n8892;
  assign n8894 = ~n8888 & n8893;
  assign n8895 = n8894 ^ x23;
  assign n9064 = n9063 ^ n8895;
  assign n8885 = n8767 ^ n8609;
  assign n8886 = ~n8768 & ~n8885;
  assign n8887 = n8886 ^ n8609;
  assign n9065 = n9064 ^ n8887;
  assign n8877 = n1404 & n5117;
  assign n8878 = x104 & n1408;
  assign n8879 = x103 & n1514;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = x105 & n1517;
  assign n8882 = n8880 & ~n8881;
  assign n8883 = ~n8877 & n8882;
  assign n8884 = n8883 ^ x20;
  assign n9066 = n9065 ^ n8884;
  assign n8874 = n8769 ^ n8598;
  assign n8875 = n8770 & n8874;
  assign n8876 = n8875 ^ n8598;
  assign n9067 = n9066 ^ n8876;
  assign n8866 = n1098 & n5792;
  assign n8867 = x106 & n1198;
  assign n8868 = x107 & n1102;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = x108 & n1201;
  assign n8871 = n8869 & ~n8870;
  assign n8872 = ~n8866 & n8871;
  assign n8873 = n8872 ^ x17;
  assign n9068 = n9067 ^ n8873;
  assign n8863 = n8771 ^ n8587;
  assign n8864 = ~n8772 & ~n8863;
  assign n8865 = n8864 ^ n8587;
  assign n9069 = n9068 ^ n8865;
  assign n8855 = n821 & n6478;
  assign n8856 = x109 & n898;
  assign n8857 = x111 & n901;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = x110 & n824;
  assign n8860 = n8858 & ~n8859;
  assign n8861 = ~n8855 & n8860;
  assign n8862 = n8861 ^ x14;
  assign n9070 = n9069 ^ n8862;
  assign n8852 = n8773 ^ n8576;
  assign n8853 = n8774 & n8852;
  assign n8854 = n8853 ^ n8576;
  assign n9071 = n9070 ^ n8854;
  assign n8844 = n596 & n7220;
  assign n8845 = x112 & n673;
  assign n8846 = x114 & n676;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = x113 & n601;
  assign n8849 = n8847 & ~n8848;
  assign n8850 = ~n8844 & n8849;
  assign n8851 = n8850 ^ x11;
  assign n9072 = n9071 ^ n8851;
  assign n8841 = n8775 ^ n8565;
  assign n8842 = ~n8776 & ~n8841;
  assign n8843 = n8842 ^ n8565;
  assign n9073 = n9072 ^ n8843;
  assign n8833 = n399 & n7987;
  assign n8834 = x115 & n478;
  assign n8835 = x116 & n402;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = x117 & n470;
  assign n8838 = n8836 & ~n8837;
  assign n8839 = ~n8833 & n8838;
  assign n8840 = n8839 ^ x8;
  assign n9074 = n9073 ^ n8840;
  assign n8830 = n8777 ^ n8554;
  assign n8831 = n8778 & n8830;
  assign n8832 = n8831 ^ n8554;
  assign n9075 = n9074 ^ n8832;
  assign n8820 = n7970 ^ x120;
  assign n8821 = n239 & n8820;
  assign n8822 = x118 & n249;
  assign n8823 = x119 & n242;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = x120 & n280;
  assign n8826 = n8824 & ~n8825;
  assign n8827 = ~n8821 & n8826;
  assign n8828 = n8827 ^ x5;
  assign n8805 = ~x122 & ~n8527;
  assign n8806 = x122 & ~n8525;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = n169 & ~n8807;
  assign n8809 = n8808 ^ x1;
  assign n8810 = n8809 ^ x123;
  assign n8803 = x122 ^ x2;
  assign n8804 = x1 & n8803;
  assign n8811 = n8810 ^ n8804;
  assign n8812 = n8811 ^ n8810;
  assign n8813 = ~x121 & n197;
  assign n8814 = n8813 ^ n8810;
  assign n8815 = n8814 ^ n8810;
  assign n8816 = ~n8812 & ~n8815;
  assign n8817 = n8816 ^ n8810;
  assign n8818 = ~x0 & ~n8817;
  assign n8819 = n8818 ^ n8810;
  assign n8829 = n8828 ^ n8819;
  assign n9076 = n9075 ^ n8829;
  assign n8783 = n8541 & ~n8550;
  assign n8784 = ~n8779 & n8783;
  assign n8785 = ~n8522 & n8784;
  assign n8786 = ~n8541 & n8550;
  assign n8787 = n8779 & n8786;
  assign n8788 = n8522 & n8787;
  assign n8789 = ~n8785 & ~n8788;
  assign n8790 = n8779 ^ n8541;
  assign n8791 = n8551 & ~n8790;
  assign n8792 = n8791 ^ n8779;
  assign n8793 = n8522 & n8792;
  assign n8794 = ~n8787 & ~n8793;
  assign n8795 = n8794 ^ n8519;
  assign n8796 = n8795 ^ n8794;
  assign n8797 = n8522 & ~n8784;
  assign n8798 = ~n8792 & ~n8797;
  assign n8799 = n8798 ^ n8794;
  assign n8800 = n8796 & ~n8799;
  assign n8801 = n8800 ^ n8794;
  assign n8802 = n8789 & n8801;
  assign n9077 = n9076 ^ n8802;
  assign n9350 = ~n8788 & n9076;
  assign n9351 = ~n8798 & ~n9350;
  assign n9352 = n8519 & ~n9351;
  assign n9353 = n8794 & n9076;
  assign n9354 = ~n8785 & ~n9353;
  assign n9355 = ~n9352 & n9354;
  assign n9306 = n458 & n8171;
  assign n9307 = x69 & n8174;
  assign n9308 = x68 & n8181;
  assign n9309 = ~n9307 & ~n9308;
  assign n9310 = x70 & n8732;
  assign n9311 = n9309 & ~n9310;
  assign n9312 = ~n9306 & n9311;
  assign n9313 = n9312 ^ x56;
  assign n9294 = x59 & n8999;
  assign n9295 = n9018 & n9294;
  assign n9296 = x60 ^ x59;
  assign n9297 = x64 & n9296;
  assign n9298 = ~n9295 & ~n9297;
  assign n9286 = n168 & n9001;
  assign n9287 = n9286 ^ x67;
  assign n9288 = n8427 & n9287;
  assign n9289 = x66 & n9005;
  assign n9290 = x65 & n9012;
  assign n9291 = ~n9289 & ~n9290;
  assign n9292 = ~n9288 & n9291;
  assign n9293 = n9292 ^ x59;
  assign n9299 = n9298 ^ n9293;
  assign n9300 = n9018 ^ x60;
  assign n9301 = x64 & n9294;
  assign n9302 = n9300 & n9301;
  assign n9303 = ~n9293 & n9302;
  assign n9304 = ~n9299 & n9303;
  assign n9305 = n9304 ^ n9299;
  assign n9314 = n9313 ^ n9305;
  assign n9283 = n9019 ^ n8991;
  assign n9284 = ~n9020 & ~n9283;
  assign n9285 = n9284 ^ n8994;
  assign n9315 = n9314 ^ n9285;
  assign n9275 = ~n653 & n7395;
  assign n9276 = x72 & n7400;
  assign n9277 = x71 & n7650;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = x73 & n7652;
  assign n9280 = n9278 & ~n9279;
  assign n9281 = ~n9275 & n9280;
  assign n9282 = n9281 ^ x53;
  assign n9316 = n9315 ^ n9282;
  assign n9272 = n9021 ^ n8975;
  assign n9273 = n9022 & n9272;
  assign n9274 = n9273 ^ n8975;
  assign n9317 = n9316 ^ n9274;
  assign n9264 = n870 & n6626;
  assign n9265 = x74 & n6884;
  assign n9266 = x76 & n6888;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = x75 & n6630;
  assign n9269 = n9267 & ~n9268;
  assign n9270 = ~n9264 & n9269;
  assign n9271 = n9270 ^ x50;
  assign n9318 = n9317 ^ n9271;
  assign n9261 = n9034 ^ n9023;
  assign n9262 = ~n9035 & ~n9261;
  assign n9263 = n9262 ^ n9026;
  assign n9319 = n9318 ^ n9263;
  assign n9253 = n1149 & n5942;
  assign n9254 = x77 & n6186;
  assign n9255 = x78 & n5947;
  assign n9256 = ~n9254 & ~n9255;
  assign n9257 = x79 & n6406;
  assign n9258 = n9256 & ~n9257;
  assign n9259 = ~n9253 & n9258;
  assign n9260 = n9259 ^ x47;
  assign n9320 = n9319 ^ n9260;
  assign n9250 = n9047 ^ n9036;
  assign n9251 = ~n9048 & n9250;
  assign n9252 = n9251 ^ n9039;
  assign n9321 = n9320 ^ n9252;
  assign n9242 = n1454 & n5262;
  assign n9243 = x80 & n5488;
  assign n9244 = x81 & n5266;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = x82 & n5491;
  assign n9247 = n9245 & ~n9246;
  assign n9248 = ~n9242 & n9247;
  assign n9249 = n9248 ^ x44;
  assign n9322 = n9321 ^ n9249;
  assign n9239 = n9049 ^ n8964;
  assign n9240 = ~n9050 & ~n9239;
  assign n9241 = n9240 ^ n8964;
  assign n9323 = n9322 ^ n9241;
  assign n9231 = n1801 & n4643;
  assign n9232 = x83 & n4653;
  assign n9233 = x85 & n5046;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = x84 & n4646;
  assign n9236 = n9234 & ~n9235;
  assign n9237 = ~n9231 & n9236;
  assign n9238 = n9237 ^ x41;
  assign n9324 = n9323 ^ n9238;
  assign n9228 = n9051 ^ n8953;
  assign n9229 = n9052 & n9228;
  assign n9230 = n9229 ^ n8953;
  assign n9325 = n9324 ^ n9230;
  assign n9220 = n2176 & n4040;
  assign n9221 = x86 & n4267;
  assign n9222 = x88 & n4270;
  assign n9223 = ~n9221 & ~n9222;
  assign n9224 = x87 & n4044;
  assign n9225 = n9223 & ~n9224;
  assign n9226 = ~n9220 & n9225;
  assign n9227 = n9226 ^ x38;
  assign n9326 = n9325 ^ n9227;
  assign n9217 = n9053 ^ n8942;
  assign n9218 = ~n9054 & ~n9217;
  assign n9219 = n9218 ^ n8942;
  assign n9327 = n9326 ^ n9219;
  assign n9209 = n2607 & n3522;
  assign n9210 = x89 & n3699;
  assign n9211 = x90 & n3526;
  assign n9212 = ~n9210 & ~n9211;
  assign n9213 = x91 & n3701;
  assign n9214 = n9212 & ~n9213;
  assign n9215 = ~n9209 & n9214;
  assign n9216 = n9215 ^ x35;
  assign n9328 = n9327 ^ n9216;
  assign n9206 = n9055 ^ n8931;
  assign n9207 = n9056 & n9206;
  assign n9208 = n9207 ^ n8931;
  assign n9329 = n9328 ^ n9208;
  assign n9198 = n3009 & n3078;
  assign n9199 = x92 & n3181;
  assign n9200 = x93 & n3013;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = x94 & n3183;
  assign n9203 = n9201 & ~n9202;
  assign n9204 = ~n9198 & n9203;
  assign n9205 = n9204 ^ x32;
  assign n9330 = n9329 ^ n9205;
  assign n9195 = n9057 ^ n8920;
  assign n9196 = ~n9058 & ~n9195;
  assign n9197 = n9196 ^ n8920;
  assign n9331 = n9330 ^ n9197;
  assign n9187 = n2527 & n3585;
  assign n9188 = x95 & n2690;
  assign n9189 = x96 & n2530;
  assign n9190 = ~n9188 & ~n9189;
  assign n9191 = x97 & n2693;
  assign n9192 = n9190 & ~n9191;
  assign n9193 = ~n9187 & n9192;
  assign n9194 = n9193 ^ x29;
  assign n9332 = n9331 ^ n9194;
  assign n9184 = n8917 ^ n8909;
  assign n9185 = ~n9060 & ~n9184;
  assign n9186 = n9185 ^ n9059;
  assign n9333 = n9332 ^ n9186;
  assign n9176 = n2102 & n4141;
  assign n9177 = x98 & n2112;
  assign n9178 = x99 & n2105;
  assign n9179 = ~n9177 & ~n9178;
  assign n9180 = x100 & n2381;
  assign n9181 = n9179 & ~n9180;
  assign n9182 = ~n9176 & n9181;
  assign n9183 = n9182 ^ x26;
  assign n9334 = n9333 ^ n9183;
  assign n9173 = n9061 ^ n8898;
  assign n9174 = n9062 & n9173;
  assign n9175 = n9174 ^ n8898;
  assign n9335 = n9334 ^ n9175;
  assign n9165 = n1746 & n4718;
  assign n9166 = x101 & n1871;
  assign n9167 = x102 & n1750;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = x103 & n1873;
  assign n9170 = n9168 & ~n9169;
  assign n9171 = ~n9165 & n9170;
  assign n9172 = n9171 ^ x23;
  assign n9336 = n9335 ^ n9172;
  assign n9162 = n9063 ^ n8887;
  assign n9163 = ~n9064 & ~n9162;
  assign n9164 = n9163 ^ n8887;
  assign n9337 = n9336 ^ n9164;
  assign n9154 = n1404 & n5351;
  assign n9155 = x104 & n1514;
  assign n9156 = x105 & n1408;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = x106 & n1517;
  assign n9159 = n9157 & ~n9158;
  assign n9160 = ~n9154 & n9159;
  assign n9161 = n9160 ^ x20;
  assign n9338 = n9337 ^ n9161;
  assign n9151 = n9065 ^ n8876;
  assign n9152 = n9066 & n9151;
  assign n9153 = n9152 ^ n8876;
  assign n9339 = n9338 ^ n9153;
  assign n9143 = n1098 & n6026;
  assign n9144 = x107 & n1198;
  assign n9145 = x108 & n1102;
  assign n9146 = ~n9144 & ~n9145;
  assign n9147 = x109 & n1201;
  assign n9148 = n9146 & ~n9147;
  assign n9149 = ~n9143 & n9148;
  assign n9150 = n9149 ^ x17;
  assign n9340 = n9339 ^ n9150;
  assign n9140 = n9067 ^ n8865;
  assign n9141 = ~n9068 & ~n9140;
  assign n9142 = n9141 ^ n8865;
  assign n9341 = n9340 ^ n9142;
  assign n9132 = n821 & n6728;
  assign n9133 = x110 & n898;
  assign n9134 = x111 & n824;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = x112 & n901;
  assign n9137 = n9135 & ~n9136;
  assign n9138 = ~n9132 & n9137;
  assign n9139 = n9138 ^ x14;
  assign n9342 = n9341 ^ n9139;
  assign n9129 = n9069 ^ n8854;
  assign n9130 = n9070 & n9129;
  assign n9131 = n9130 ^ n8854;
  assign n9343 = n9342 ^ n9131;
  assign n9121 = n596 & n7481;
  assign n9122 = x113 & n673;
  assign n9123 = x114 & n601;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = x115 & n676;
  assign n9126 = n9124 & ~n9125;
  assign n9127 = ~n9121 & n9126;
  assign n9128 = n9127 ^ x11;
  assign n9344 = n9343 ^ n9128;
  assign n9118 = n9071 ^ n8843;
  assign n9119 = ~n9072 & ~n9118;
  assign n9120 = n9119 ^ n8843;
  assign n9345 = n9344 ^ n9120;
  assign n9110 = n399 & n8265;
  assign n9111 = x116 & n478;
  assign n9112 = x117 & n402;
  assign n9113 = ~n9111 & ~n9112;
  assign n9114 = x118 & n470;
  assign n9115 = n9113 & ~n9114;
  assign n9116 = ~n9110 & n9115;
  assign n9117 = n9116 ^ x8;
  assign n9346 = n9345 ^ n9117;
  assign n9107 = n9073 ^ n8832;
  assign n9108 = n9074 & n9107;
  assign n9109 = n9108 ^ n8832;
  assign n9347 = n9346 ^ n9109;
  assign n9104 = n9075 ^ n8819;
  assign n9105 = n8829 & ~n9104;
  assign n9106 = n9105 ^ n9075;
  assign n9348 = n9347 ^ n9106;
  assign n9094 = n8249 ^ x121;
  assign n9095 = n239 & n9094;
  assign n9096 = x119 & n249;
  assign n9097 = x121 & n280;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = x120 & n242;
  assign n9100 = n9098 & ~n9099;
  assign n9101 = ~n9095 & n9100;
  assign n9102 = n9101 ^ x5;
  assign n9080 = x123 ^ x122;
  assign n9081 = ~n8807 & n9080;
  assign n9082 = n169 & ~n9081;
  assign n9083 = n9082 ^ x1;
  assign n9084 = n9083 ^ x124;
  assign n9078 = x1 & x123;
  assign n9079 = n9078 ^ x2;
  assign n9085 = n9084 ^ n9079;
  assign n9086 = n9085 ^ n9084;
  assign n9087 = x122 & n197;
  assign n9088 = n9087 ^ n9084;
  assign n9089 = n9088 ^ n9084;
  assign n9090 = n9086 & ~n9089;
  assign n9091 = n9090 ^ n9084;
  assign n9092 = ~x0 & n9091;
  assign n9093 = n9092 ^ n9084;
  assign n9103 = n9102 ^ n9093;
  assign n9349 = n9348 ^ n9103;
  assign n9356 = n9355 ^ n9349;
  assign n9628 = ~n9106 & ~n9347;
  assign n9629 = n9093 & ~n9102;
  assign n9630 = n9628 & n9629;
  assign n9631 = n9106 & n9347;
  assign n9632 = ~n9093 & n9102;
  assign n9633 = n9631 & n9632;
  assign n9634 = ~n9630 & ~n9633;
  assign n9639 = n9628 ^ n9093;
  assign n9640 = n9106 ^ n9102;
  assign n9641 = n9640 ^ n9347;
  assign n9642 = n9631 & n9641;
  assign n9643 = n9642 ^ n9641;
  assign n9644 = n9639 & ~n9643;
  assign n9645 = n9644 ^ n9093;
  assign n9635 = n9631 ^ n9093;
  assign n9636 = ~n9103 & ~n9635;
  assign n9637 = n9636 ^ n9093;
  assign n9638 = ~n9628 & ~n9637;
  assign n9646 = n9645 ^ n9638;
  assign n9647 = ~n9355 & n9646;
  assign n9648 = n9647 ^ n9638;
  assign n9649 = n9634 & ~n9648;
  assign n9590 = n956 & n6626;
  assign n9591 = x75 & n6884;
  assign n9592 = x76 & n6630;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = x77 & n6888;
  assign n9595 = n9593 & ~n9594;
  assign n9596 = ~n9590 & n9595;
  assign n9597 = n9596 ^ x50;
  assign n9587 = n9317 ^ n9263;
  assign n9588 = n9318 & n9587;
  assign n9589 = n9588 ^ n9263;
  assign n9598 = n9597 ^ n9589;
  assign n9575 = n517 & n8171;
  assign n9576 = x70 & n8174;
  assign n9577 = x69 & n8181;
  assign n9578 = ~n9576 & ~n9577;
  assign n9579 = x71 & n8732;
  assign n9580 = n9578 & ~n9579;
  assign n9581 = ~n9575 & n9580;
  assign n9582 = n9581 ^ x56;
  assign n9572 = ~n9293 & ~n9298;
  assign n9567 = x65 ^ x60;
  assign n9568 = n9296 & ~n9567;
  assign n9569 = n9568 ^ x59;
  assign n9570 = n9569 ^ x61;
  assign n9564 = x59 & x60;
  assign n9565 = n9564 ^ x61;
  assign n9566 = ~x64 & n9565;
  assign n9571 = n9570 ^ n9566;
  assign n9573 = n9572 ^ n9571;
  assign n9555 = n321 & n9002;
  assign n9556 = x66 & n9012;
  assign n9557 = n8427 & ~n9001;
  assign n9558 = x68 & n9557;
  assign n9559 = ~n9556 & ~n9558;
  assign n9560 = x67 & n9005;
  assign n9561 = n9559 & ~n9560;
  assign n9562 = ~n9555 & n9561;
  assign n9563 = n9562 ^ x59;
  assign n9574 = n9573 ^ n9563;
  assign n9583 = n9582 ^ n9574;
  assign n9552 = n9305 ^ n9285;
  assign n9553 = n9314 & n9552;
  assign n9554 = n9553 ^ n9285;
  assign n9584 = n9583 ^ n9554;
  assign n9544 = ~n721 & n7395;
  assign n9545 = x72 & n7650;
  assign n9546 = x73 & n7400;
  assign n9547 = ~n9545 & ~n9546;
  assign n9548 = x74 & n7652;
  assign n9549 = n9547 & ~n9548;
  assign n9550 = ~n9544 & n9549;
  assign n9551 = n9550 ^ x53;
  assign n9585 = n9584 ^ n9551;
  assign n9541 = n9315 ^ n9274;
  assign n9542 = ~n9316 & ~n9541;
  assign n9543 = n9542 ^ n9274;
  assign n9586 = n9585 ^ n9543;
  assign n9599 = n9598 ^ n9586;
  assign n9533 = n1242 & n5942;
  assign n9534 = x78 & n6186;
  assign n9535 = x79 & n5947;
  assign n9536 = ~n9534 & ~n9535;
  assign n9537 = x80 & n6406;
  assign n9538 = n9536 & ~n9537;
  assign n9539 = ~n9533 & n9538;
  assign n9540 = n9539 ^ x47;
  assign n9600 = n9599 ^ n9540;
  assign n9530 = n9319 ^ n9252;
  assign n9531 = ~n9320 & ~n9530;
  assign n9532 = n9531 ^ n9252;
  assign n9601 = n9600 ^ n9532;
  assign n9522 = n1560 & n5262;
  assign n9523 = x81 & n5488;
  assign n9524 = x82 & n5266;
  assign n9525 = ~n9523 & ~n9524;
  assign n9526 = x83 & n5491;
  assign n9527 = n9525 & ~n9526;
  assign n9528 = ~n9522 & n9527;
  assign n9529 = n9528 ^ x44;
  assign n9602 = n9601 ^ n9529;
  assign n9519 = n9321 ^ n9241;
  assign n9520 = n9322 & n9519;
  assign n9521 = n9520 ^ n9241;
  assign n9603 = n9602 ^ n9521;
  assign n9511 = n1920 & n4643;
  assign n9512 = x84 & n4653;
  assign n9513 = x86 & n5046;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = x85 & n4646;
  assign n9516 = n9514 & ~n9515;
  assign n9517 = ~n9511 & n9516;
  assign n9518 = n9517 ^ x41;
  assign n9604 = n9603 ^ n9518;
  assign n9508 = n9323 ^ n9230;
  assign n9509 = ~n9324 & ~n9508;
  assign n9510 = n9509 ^ n9230;
  assign n9605 = n9604 ^ n9510;
  assign n9500 = n2310 & n4040;
  assign n9501 = x87 & n4267;
  assign n9502 = x89 & n4270;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = x88 & n4044;
  assign n9505 = n9503 & ~n9504;
  assign n9506 = ~n9500 & n9505;
  assign n9507 = n9506 ^ x38;
  assign n9606 = n9605 ^ n9507;
  assign n9497 = n9325 ^ n9219;
  assign n9498 = n9326 & n9497;
  assign n9499 = n9498 ^ n9219;
  assign n9607 = n9606 ^ n9499;
  assign n9489 = n2755 & n3522;
  assign n9490 = x90 & n3699;
  assign n9491 = x91 & n3526;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = x92 & n3701;
  assign n9494 = n9492 & ~n9493;
  assign n9495 = ~n9489 & n9494;
  assign n9496 = n9495 ^ x35;
  assign n9608 = n9607 ^ n9496;
  assign n9486 = n9327 ^ n9208;
  assign n9487 = ~n9328 & ~n9486;
  assign n9488 = n9487 ^ n9208;
  assign n9609 = n9608 ^ n9488;
  assign n9478 = n3009 & n3247;
  assign n9479 = x93 & n3181;
  assign n9480 = x94 & n3013;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = x95 & n3183;
  assign n9483 = n9481 & ~n9482;
  assign n9484 = ~n9478 & n9483;
  assign n9485 = n9484 ^ x32;
  assign n9610 = n9609 ^ n9485;
  assign n9475 = n9329 ^ n9197;
  assign n9476 = n9330 & n9475;
  assign n9477 = n9476 ^ n9197;
  assign n9611 = n9610 ^ n9477;
  assign n9467 = n2527 & n3763;
  assign n9468 = x96 & n2690;
  assign n9469 = x97 & n2530;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = x98 & n2693;
  assign n9472 = n9470 & ~n9471;
  assign n9473 = ~n9467 & n9472;
  assign n9474 = n9473 ^ x29;
  assign n9612 = n9611 ^ n9474;
  assign n9464 = n9194 ^ n9186;
  assign n9465 = n9332 & n9464;
  assign n9466 = n9465 ^ n9331;
  assign n9613 = n9612 ^ n9466;
  assign n9456 = n2102 & n4323;
  assign n9457 = x99 & n2112;
  assign n9458 = x100 & n2105;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = x101 & n2381;
  assign n9461 = n9459 & ~n9460;
  assign n9462 = ~n9456 & n9461;
  assign n9463 = n9462 ^ x26;
  assign n9614 = n9613 ^ n9463;
  assign n9453 = n9333 ^ n9175;
  assign n9454 = n9334 & n9453;
  assign n9455 = n9454 ^ n9175;
  assign n9615 = n9614 ^ n9455;
  assign n9445 = n1746 & n4912;
  assign n9446 = x102 & n1871;
  assign n9447 = x103 & n1750;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = x104 & n1873;
  assign n9450 = n9448 & ~n9449;
  assign n9451 = ~n9445 & n9450;
  assign n9452 = n9451 ^ x23;
  assign n9616 = n9615 ^ n9452;
  assign n9442 = n9335 ^ n9164;
  assign n9443 = ~n9336 & ~n9442;
  assign n9444 = n9443 ^ n9164;
  assign n9617 = n9616 ^ n9444;
  assign n9434 = n1404 & n5578;
  assign n9435 = x105 & n1514;
  assign n9436 = x106 & n1408;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = x107 & n1517;
  assign n9439 = n9437 & ~n9438;
  assign n9440 = ~n9434 & n9439;
  assign n9441 = n9440 ^ x20;
  assign n9618 = n9617 ^ n9441;
  assign n9431 = n9337 ^ n9153;
  assign n9432 = n9338 & n9431;
  assign n9433 = n9432 ^ n9153;
  assign n9619 = n9618 ^ n9433;
  assign n9423 = n1098 & n6250;
  assign n9424 = x108 & n1198;
  assign n9425 = x109 & n1102;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = x110 & n1201;
  assign n9428 = n9426 & ~n9427;
  assign n9429 = ~n9423 & n9428;
  assign n9430 = n9429 ^ x17;
  assign n9620 = n9619 ^ n9430;
  assign n9420 = n9339 ^ n9142;
  assign n9421 = ~n9340 & ~n9420;
  assign n9422 = n9421 ^ n9142;
  assign n9621 = n9620 ^ n9422;
  assign n9412 = n821 & n6975;
  assign n9413 = x111 & n898;
  assign n9414 = x112 & n824;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = x113 & n901;
  assign n9417 = n9415 & ~n9416;
  assign n9418 = ~n9412 & n9417;
  assign n9419 = n9418 ^ x14;
  assign n9622 = n9621 ^ n9419;
  assign n9409 = n9341 ^ n9131;
  assign n9410 = n9342 & n9409;
  assign n9411 = n9410 ^ n9131;
  assign n9623 = n9622 ^ n9411;
  assign n9401 = n596 & n7730;
  assign n9402 = x114 & n673;
  assign n9403 = x116 & n676;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = x115 & n601;
  assign n9406 = n9404 & ~n9405;
  assign n9407 = ~n9401 & n9406;
  assign n9408 = n9407 ^ x11;
  assign n9624 = n9623 ^ n9408;
  assign n9398 = n9343 ^ n9120;
  assign n9399 = ~n9344 & ~n9398;
  assign n9400 = n9399 ^ n9120;
  assign n9625 = n9624 ^ n9400;
  assign n9387 = n8528 ^ x122;
  assign n9388 = n239 & n9387;
  assign n9389 = x120 & n249;
  assign n9390 = x121 & n242;
  assign n9391 = ~n9389 & ~n9390;
  assign n9392 = x122 & n280;
  assign n9393 = n9391 & ~n9392;
  assign n9394 = ~n9388 & n9393;
  assign n9395 = n9394 ^ x5;
  assign n9379 = n399 & n8542;
  assign n9380 = x117 & n478;
  assign n9381 = x119 & n470;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = x118 & n402;
  assign n9384 = n9382 & ~n9383;
  assign n9385 = ~n9379 & n9384;
  assign n9386 = n9385 ^ x8;
  assign n9396 = n9395 ^ n9386;
  assign n9362 = x124 & n8806;
  assign n9363 = ~x123 & ~n9362;
  assign n9364 = ~x124 & n8805;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = n9365 ^ x124;
  assign n9367 = n169 & ~n9366;
  assign n9368 = n9367 ^ x1;
  assign n9369 = n9368 ^ x125;
  assign n9360 = x124 ^ x2;
  assign n9361 = x1 & n9360;
  assign n9370 = n9369 ^ n9361;
  assign n9371 = n9370 ^ n9369;
  assign n9372 = ~x123 & n197;
  assign n9373 = n9372 ^ n9369;
  assign n9374 = n9373 ^ n9369;
  assign n9375 = ~n9371 & ~n9374;
  assign n9376 = n9375 ^ n9369;
  assign n9377 = ~x0 & ~n9376;
  assign n9378 = n9377 ^ n9369;
  assign n9397 = n9396 ^ n9378;
  assign n9626 = n9625 ^ n9397;
  assign n9357 = n9345 ^ n9109;
  assign n9358 = n9346 & n9357;
  assign n9359 = n9358 ^ n9109;
  assign n9627 = n9626 ^ n9359;
  assign n9650 = n9649 ^ n9627;
  assign n9951 = ~n9627 & ~n9628;
  assign n9952 = n9629 & ~n9951;
  assign n9953 = n9355 & ~n9952;
  assign n9954 = n9627 & ~n9633;
  assign n9955 = ~n9645 & ~n9954;
  assign n9956 = ~n9953 & ~n9955;
  assign n9957 = n9632 ^ n9106;
  assign n9958 = n9348 & n9957;
  assign n9959 = n9958 ^ n9106;
  assign n9960 = n9627 & ~n9959;
  assign n9961 = ~n9956 & ~n9960;
  assign n9910 = n789 & n7395;
  assign n9911 = x74 & n7400;
  assign n9912 = x73 & n7650;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = x75 & n7652;
  assign n9915 = n9913 & ~n9914;
  assign n9916 = ~n9910 & n9915;
  assign n9917 = n9916 ^ x53;
  assign n9907 = n9584 ^ n9543;
  assign n9908 = n9585 & n9907;
  assign n9909 = n9908 ^ n9543;
  assign n9918 = n9917 ^ n9909;
  assign n9896 = n420 & n9002;
  assign n9897 = x67 & n9012;
  assign n9898 = x69 & n9557;
  assign n9899 = ~n9897 & ~n9898;
  assign n9900 = x68 & n9005;
  assign n9901 = n9899 & ~n9900;
  assign n9902 = ~n9896 & n9901;
  assign n9877 = x62 ^ x61;
  assign n9878 = n9296 & n9877;
  assign n9879 = n142 & n9878;
  assign n9880 = x61 & ~n9296;
  assign n9881 = n9880 ^ n9564;
  assign n9882 = ~n9879 & ~n9881;
  assign n9883 = x65 & ~n9882;
  assign n9884 = n9564 ^ x62;
  assign n9885 = n9884 ^ n9564;
  assign n9886 = ~n9296 & n9885;
  assign n9887 = n9886 ^ n9564;
  assign n9888 = n9877 & n9887;
  assign n9889 = x64 & n9888;
  assign n9890 = n152 & n9877;
  assign n9891 = x66 & n9296;
  assign n9892 = ~n9890 & n9891;
  assign n9893 = ~n9889 & ~n9892;
  assign n9894 = ~n9883 & n9893;
  assign n9871 = x61 ^ x59;
  assign n9872 = x64 & n9871;
  assign n9873 = n9872 ^ n233;
  assign n9874 = ~n9296 & ~n9873;
  assign n9875 = n9874 ^ n233;
  assign n9876 = x62 & ~n9875;
  assign n9895 = n9894 ^ n9876;
  assign n9903 = n9902 ^ n9895;
  assign n9867 = n9571 ^ x59;
  assign n9868 = n9867 ^ n9562;
  assign n9869 = ~n9573 & ~n9868;
  assign n9870 = n9869 ^ n9562;
  assign n9904 = n9903 ^ n9870;
  assign n9859 = n575 & n8171;
  assign n9860 = x71 & n8174;
  assign n9861 = x70 & n8181;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = x72 & n8732;
  assign n9864 = n9862 & ~n9863;
  assign n9865 = ~n9859 & n9864;
  assign n9866 = n9865 ^ x56;
  assign n9905 = n9904 ^ n9866;
  assign n9856 = n9582 ^ n9554;
  assign n9857 = ~n9583 & ~n9856;
  assign n9858 = n9857 ^ n9554;
  assign n9906 = n9905 ^ n9858;
  assign n9919 = n9918 ^ n9906;
  assign n9847 = n1340 & n5942;
  assign n9848 = x79 & n6186;
  assign n9849 = x81 & n6406;
  assign n9850 = ~n9848 & ~n9849;
  assign n9851 = x80 & n5947;
  assign n9852 = n9850 & ~n9851;
  assign n9853 = ~n9847 & n9852;
  assign n9854 = n9853 ^ x47;
  assign n9839 = n1041 & n6626;
  assign n9840 = x77 & n6630;
  assign n9841 = x76 & n6884;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = x78 & n6888;
  assign n9844 = n9842 & ~n9843;
  assign n9845 = ~n9839 & n9844;
  assign n9846 = n9845 ^ x50;
  assign n9855 = n9854 ^ n9846;
  assign n9920 = n9919 ^ n9855;
  assign n9836 = n9597 ^ n9586;
  assign n9837 = ~n9598 & ~n9836;
  assign n9838 = n9837 ^ n9589;
  assign n9921 = n9920 ^ n9838;
  assign n9833 = n9599 ^ n9532;
  assign n9834 = n9600 & n9833;
  assign n9835 = n9834 ^ n9532;
  assign n9922 = n9921 ^ n9835;
  assign n9825 = n1667 & n5262;
  assign n9826 = x82 & n5488;
  assign n9827 = x84 & n5491;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = x83 & n5266;
  assign n9830 = n9828 & ~n9829;
  assign n9831 = ~n9825 & n9830;
  assign n9832 = n9831 ^ x44;
  assign n9923 = n9922 ^ n9832;
  assign n9822 = n9601 ^ n9521;
  assign n9823 = ~n9602 & ~n9822;
  assign n9824 = n9823 ^ n9521;
  assign n9924 = n9923 ^ n9824;
  assign n9814 = n2039 & n4643;
  assign n9815 = x85 & n4653;
  assign n9816 = x86 & n4646;
  assign n9817 = ~n9815 & ~n9816;
  assign n9818 = x87 & n5046;
  assign n9819 = n9817 & ~n9818;
  assign n9820 = ~n9814 & n9819;
  assign n9821 = n9820 ^ x41;
  assign n9925 = n9924 ^ n9821;
  assign n9811 = n9603 ^ n9510;
  assign n9812 = n9604 & n9811;
  assign n9813 = n9812 ^ n9510;
  assign n9926 = n9925 ^ n9813;
  assign n9803 = n2448 & n4040;
  assign n9804 = x88 & n4267;
  assign n9805 = x90 & n4270;
  assign n9806 = ~n9804 & ~n9805;
  assign n9807 = x89 & n4044;
  assign n9808 = n9806 & ~n9807;
  assign n9809 = ~n9803 & n9808;
  assign n9810 = n9809 ^ x38;
  assign n9927 = n9926 ^ n9810;
  assign n9800 = n9605 ^ n9499;
  assign n9801 = ~n9606 & ~n9800;
  assign n9802 = n9801 ^ n9499;
  assign n9928 = n9927 ^ n9802;
  assign n9792 = n2901 & n3522;
  assign n9793 = x91 & n3699;
  assign n9794 = x93 & n3701;
  assign n9795 = ~n9793 & ~n9794;
  assign n9796 = x92 & n3526;
  assign n9797 = n9795 & ~n9796;
  assign n9798 = ~n9792 & n9797;
  assign n9799 = n9798 ^ x35;
  assign n9929 = n9928 ^ n9799;
  assign n9789 = n9607 ^ n9488;
  assign n9790 = n9608 & n9789;
  assign n9791 = n9790 ^ n9488;
  assign n9930 = n9929 ^ n9791;
  assign n9781 = n3009 & n3403;
  assign n9782 = x94 & n3181;
  assign n9783 = x95 & n3013;
  assign n9784 = ~n9782 & ~n9783;
  assign n9785 = x96 & n3183;
  assign n9786 = n9784 & ~n9785;
  assign n9787 = ~n9781 & n9786;
  assign n9788 = n9787 ^ x32;
  assign n9931 = n9930 ^ n9788;
  assign n9778 = n9609 ^ n9477;
  assign n9779 = ~n9610 & ~n9778;
  assign n9780 = n9779 ^ n9477;
  assign n9932 = n9931 ^ n9780;
  assign n9770 = n2527 & n3943;
  assign n9771 = x97 & n2690;
  assign n9772 = x98 & n2530;
  assign n9773 = ~n9771 & ~n9772;
  assign n9774 = x99 & n2693;
  assign n9775 = n9773 & ~n9774;
  assign n9776 = ~n9770 & n9775;
  assign n9777 = n9776 ^ x29;
  assign n9933 = n9932 ^ n9777;
  assign n9767 = n9474 ^ n9466;
  assign n9768 = ~n9612 & ~n9767;
  assign n9769 = n9768 ^ n9611;
  assign n9934 = n9933 ^ n9769;
  assign n9759 = n2102 & n4509;
  assign n9760 = x100 & n2112;
  assign n9761 = x102 & n2381;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = x101 & n2105;
  assign n9764 = n9762 & ~n9763;
  assign n9765 = ~n9759 & n9764;
  assign n9766 = n9765 ^ x26;
  assign n9935 = n9934 ^ n9766;
  assign n9756 = n9613 ^ n9455;
  assign n9757 = n9614 & n9756;
  assign n9758 = n9757 ^ n9455;
  assign n9936 = n9935 ^ n9758;
  assign n9748 = n1746 & n5117;
  assign n9749 = x103 & n1871;
  assign n9750 = x104 & n1750;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = x105 & n1873;
  assign n9753 = n9751 & ~n9752;
  assign n9754 = ~n9748 & n9753;
  assign n9755 = n9754 ^ x23;
  assign n9937 = n9936 ^ n9755;
  assign n9745 = n9615 ^ n9444;
  assign n9746 = ~n9616 & ~n9745;
  assign n9747 = n9746 ^ n9444;
  assign n9938 = n9937 ^ n9747;
  assign n9737 = n1404 & n5792;
  assign n9738 = x106 & n1514;
  assign n9739 = x107 & n1408;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = x108 & n1517;
  assign n9742 = n9740 & ~n9741;
  assign n9743 = ~n9737 & n9742;
  assign n9744 = n9743 ^ x20;
  assign n9939 = n9938 ^ n9744;
  assign n9734 = n9617 ^ n9433;
  assign n9735 = n9618 & n9734;
  assign n9736 = n9735 ^ n9433;
  assign n9940 = n9939 ^ n9736;
  assign n9726 = n1098 & n6478;
  assign n9727 = x109 & n1198;
  assign n9728 = x110 & n1102;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = x111 & n1201;
  assign n9731 = n9729 & ~n9730;
  assign n9732 = ~n9726 & n9731;
  assign n9733 = n9732 ^ x17;
  assign n9941 = n9940 ^ n9733;
  assign n9723 = n9619 ^ n9422;
  assign n9724 = ~n9620 & ~n9723;
  assign n9725 = n9724 ^ n9422;
  assign n9942 = n9941 ^ n9725;
  assign n9715 = n821 & n7220;
  assign n9716 = x112 & n898;
  assign n9717 = x114 & n901;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = x113 & n824;
  assign n9720 = n9718 & ~n9719;
  assign n9721 = ~n9715 & n9720;
  assign n9722 = n9721 ^ x14;
  assign n9943 = n9942 ^ n9722;
  assign n9712 = n9621 ^ n9411;
  assign n9713 = n9622 & n9712;
  assign n9714 = n9713 ^ n9411;
  assign n9944 = n9943 ^ n9714;
  assign n9704 = n596 & n7987;
  assign n9705 = x115 & n673;
  assign n9706 = x117 & n676;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = x116 & n601;
  assign n9709 = n9707 & ~n9708;
  assign n9710 = ~n9704 & n9709;
  assign n9711 = n9710 ^ x11;
  assign n9945 = n9944 ^ n9711;
  assign n9701 = n9623 ^ n9400;
  assign n9702 = ~n9624 & ~n9701;
  assign n9703 = n9702 ^ n9400;
  assign n9946 = n9945 ^ n9703;
  assign n9691 = n8807 ^ x123;
  assign n9692 = n239 & n9691;
  assign n9693 = x121 & n249;
  assign n9694 = x123 & n280;
  assign n9695 = ~n9693 & ~n9694;
  assign n9696 = x122 & n242;
  assign n9697 = n9695 & ~n9696;
  assign n9698 = ~n9692 & n9697;
  assign n9699 = n9698 ^ x5;
  assign n9683 = n399 & n8820;
  assign n9684 = x118 & n478;
  assign n9685 = x119 & n402;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = x120 & n470;
  assign n9688 = n9686 & ~n9687;
  assign n9689 = ~n9683 & n9688;
  assign n9690 = n9689 ^ x8;
  assign n9700 = n9699 ^ n9690;
  assign n9947 = n9946 ^ n9700;
  assign n9672 = ~x124 & x125;
  assign n9673 = ~n9365 & n9672;
  assign n9674 = x124 & ~x125;
  assign n9675 = ~n9363 & n9674;
  assign n9676 = ~n9673 & ~n9675;
  assign n9677 = n169 & n9676;
  assign n9678 = n9677 ^ x1;
  assign n9679 = n9678 ^ x126;
  assign n9660 = x125 ^ x2;
  assign n9661 = n9660 ^ x1;
  assign n9662 = n9661 ^ n9660;
  assign n9663 = n9662 ^ x0;
  assign n9664 = n9660 ^ x125;
  assign n9665 = n9664 ^ x124;
  assign n9666 = ~x124 & ~n9665;
  assign n9667 = n9666 ^ n9660;
  assign n9668 = n9667 ^ x124;
  assign n9669 = n9663 & ~n9668;
  assign n9670 = n9669 ^ n9666;
  assign n9671 = n9670 ^ x124;
  assign n9680 = n9679 ^ n9671;
  assign n9681 = ~x0 & ~n9680;
  assign n9682 = n9681 ^ n9679;
  assign n9948 = n9947 ^ n9682;
  assign n9652 = n9625 ^ n9386;
  assign n9657 = n9625 ^ n9359;
  assign n9658 = n9652 & n9657;
  assign n9659 = n9658 ^ n9359;
  assign n9949 = n9948 ^ n9659;
  assign n9651 = n9395 ^ n9378;
  assign n9653 = n9652 ^ n9359;
  assign n9654 = n9653 ^ n9395;
  assign n9655 = ~n9651 & ~n9654;
  assign n9656 = n9655 ^ n9378;
  assign n9950 = n9949 ^ n9656;
  assign n9962 = n9961 ^ n9950;
  assign n10220 = ~n653 & n8171;
  assign n10221 = x72 & n8174;
  assign n10222 = x71 & n8181;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = x73 & n8732;
  assign n10225 = n10223 & ~n10224;
  assign n10226 = ~n10220 & n10225;
  assign n10227 = n10226 ^ x56;
  assign n10217 = n9904 ^ n9858;
  assign n10218 = ~n9905 & ~n10217;
  assign n10219 = n10218 ^ n9858;
  assign n10228 = n10227 ^ n10219;
  assign n10205 = ~n9571 & ~n9572;
  assign n10206 = n9903 ^ n9562;
  assign n10207 = ~n9563 & n10206;
  assign n10208 = ~n10205 & n10207;
  assign n10209 = n9571 & n9572;
  assign n10210 = n10209 ^ n9895;
  assign n10211 = n9902 ^ x59;
  assign n10212 = n10211 ^ n9895;
  assign n10213 = ~n10210 & ~n10212;
  assign n10214 = n10213 ^ n10209;
  assign n10215 = ~n10208 & ~n10214;
  assign n10196 = n458 & n9002;
  assign n10197 = x68 & n9012;
  assign n10198 = x70 & n9557;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = x69 & n9005;
  assign n10201 = n10199 & ~n10200;
  assign n10202 = ~n10196 & n10201;
  assign n10203 = n10202 ^ x59;
  assign n10175 = x62 & n9875;
  assign n10176 = n9894 & n10175;
  assign n10179 = n168 & n9877;
  assign n10180 = n10179 ^ x67;
  assign n10181 = n9296 & n10180;
  assign n10182 = x65 & n9888;
  assign n10183 = x66 & n9881;
  assign n10184 = ~n10182 & ~n10183;
  assign n10185 = ~n10181 & n10184;
  assign n10186 = n10185 ^ x62;
  assign n10177 = x63 ^ x62;
  assign n10178 = x64 & n10177;
  assign n10187 = n10186 ^ n10178;
  assign n10188 = n10187 ^ n10185;
  assign n10189 = n10188 ^ n10187;
  assign n10190 = n10187 ^ n10178;
  assign n10191 = n10190 ^ n10187;
  assign n10192 = n10189 & ~n10191;
  assign n10193 = n10192 ^ n10187;
  assign n10194 = n10176 & n10193;
  assign n10195 = n10194 ^ n10187;
  assign n10204 = n10203 ^ n10195;
  assign n10216 = n10215 ^ n10204;
  assign n10229 = n10228 ^ n10216;
  assign n10167 = n870 & n7395;
  assign n10168 = x74 & n7650;
  assign n10169 = x75 & n7400;
  assign n10170 = ~n10168 & ~n10169;
  assign n10171 = x76 & n7652;
  assign n10172 = n10170 & ~n10171;
  assign n10173 = ~n10167 & n10172;
  assign n10174 = n10173 ^ x53;
  assign n10230 = n10229 ^ n10174;
  assign n10164 = n9917 ^ n9906;
  assign n10165 = ~n9918 & n10164;
  assign n10166 = n10165 ^ n9909;
  assign n10231 = n10230 ^ n10166;
  assign n10160 = n9919 ^ n9838;
  assign n10161 = n9919 ^ n9846;
  assign n10162 = ~n10160 & ~n10161;
  assign n10163 = n10162 ^ n9838;
  assign n10232 = n10231 ^ n10163;
  assign n10152 = n1149 & n6626;
  assign n10153 = x77 & n6884;
  assign n10154 = x79 & n6888;
  assign n10155 = ~n10153 & ~n10154;
  assign n10156 = x78 & n6630;
  assign n10157 = n10155 & ~n10156;
  assign n10158 = ~n10152 & n10157;
  assign n10159 = n10158 ^ x50;
  assign n10233 = n10232 ^ n10159;
  assign n10144 = n1454 & n5942;
  assign n10145 = x80 & n6186;
  assign n10146 = x82 & n6406;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = x81 & n5947;
  assign n10149 = n10147 & ~n10148;
  assign n10150 = ~n10144 & n10149;
  assign n10151 = n10150 ^ x47;
  assign n10234 = n10233 ^ n10151;
  assign n10141 = n9854 ^ n9835;
  assign n10142 = n9921 & ~n10141;
  assign n10143 = n10142 ^ n9835;
  assign n10235 = n10234 ^ n10143;
  assign n10133 = n1801 & n5262;
  assign n10134 = x83 & n5488;
  assign n10135 = x84 & n5266;
  assign n10136 = ~n10134 & ~n10135;
  assign n10137 = x85 & n5491;
  assign n10138 = n10136 & ~n10137;
  assign n10139 = ~n10133 & n10138;
  assign n10140 = n10139 ^ x44;
  assign n10236 = n10235 ^ n10140;
  assign n10130 = n9922 ^ n9824;
  assign n10131 = ~n9923 & ~n10130;
  assign n10132 = n10131 ^ n9824;
  assign n10237 = n10236 ^ n10132;
  assign n10122 = n2176 & n4643;
  assign n10123 = x86 & n4653;
  assign n10124 = x88 & n5046;
  assign n10125 = ~n10123 & ~n10124;
  assign n10126 = x87 & n4646;
  assign n10127 = n10125 & ~n10126;
  assign n10128 = ~n10122 & n10127;
  assign n10129 = n10128 ^ x41;
  assign n10238 = n10237 ^ n10129;
  assign n10119 = n9924 ^ n9813;
  assign n10120 = n9925 & n10119;
  assign n10121 = n10120 ^ n9813;
  assign n10239 = n10238 ^ n10121;
  assign n10111 = n2607 & n4040;
  assign n10112 = x89 & n4267;
  assign n10113 = x91 & n4270;
  assign n10114 = ~n10112 & ~n10113;
  assign n10115 = x90 & n4044;
  assign n10116 = n10114 & ~n10115;
  assign n10117 = ~n10111 & n10116;
  assign n10118 = n10117 ^ x38;
  assign n10240 = n10239 ^ n10118;
  assign n10108 = n9926 ^ n9802;
  assign n10109 = ~n9927 & ~n10108;
  assign n10110 = n10109 ^ n9802;
  assign n10241 = n10240 ^ n10110;
  assign n10100 = n3078 & n3522;
  assign n10101 = x92 & n3699;
  assign n10102 = x94 & n3701;
  assign n10103 = ~n10101 & ~n10102;
  assign n10104 = x93 & n3526;
  assign n10105 = n10103 & ~n10104;
  assign n10106 = ~n10100 & n10105;
  assign n10107 = n10106 ^ x35;
  assign n10242 = n10241 ^ n10107;
  assign n10097 = n9928 ^ n9791;
  assign n10098 = n9929 & n10097;
  assign n10099 = n10098 ^ n9791;
  assign n10243 = n10242 ^ n10099;
  assign n10089 = n3009 & n3585;
  assign n10090 = x95 & n3181;
  assign n10091 = x96 & n3013;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = x97 & n3183;
  assign n10094 = n10092 & ~n10093;
  assign n10095 = ~n10089 & n10094;
  assign n10096 = n10095 ^ x32;
  assign n10244 = n10243 ^ n10096;
  assign n10086 = n9930 ^ n9780;
  assign n10087 = ~n9931 & ~n10086;
  assign n10088 = n10087 ^ n9780;
  assign n10245 = n10244 ^ n10088;
  assign n10078 = n2527 & n4141;
  assign n10079 = x98 & n2690;
  assign n10080 = x99 & n2530;
  assign n10081 = ~n10079 & ~n10080;
  assign n10082 = x100 & n2693;
  assign n10083 = n10081 & ~n10082;
  assign n10084 = ~n10078 & n10083;
  assign n10085 = n10084 ^ x29;
  assign n10246 = n10245 ^ n10085;
  assign n10075 = n9777 ^ n9769;
  assign n10076 = ~n9933 & n10075;
  assign n10077 = n10076 ^ n9932;
  assign n10247 = n10246 ^ n10077;
  assign n10067 = n2102 & n4718;
  assign n10068 = x101 & n2112;
  assign n10069 = x102 & n2105;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 = x103 & n2381;
  assign n10072 = n10070 & ~n10071;
  assign n10073 = ~n10067 & n10072;
  assign n10074 = n10073 ^ x26;
  assign n10248 = n10247 ^ n10074;
  assign n10064 = n9934 ^ n9758;
  assign n10065 = ~n9935 & ~n10064;
  assign n10066 = n10065 ^ n9758;
  assign n10249 = n10248 ^ n10066;
  assign n10056 = n1746 & n5351;
  assign n10057 = x105 & n1750;
  assign n10058 = x104 & n1871;
  assign n10059 = ~n10057 & ~n10058;
  assign n10060 = x106 & n1873;
  assign n10061 = n10059 & ~n10060;
  assign n10062 = ~n10056 & n10061;
  assign n10063 = n10062 ^ x23;
  assign n10250 = n10249 ^ n10063;
  assign n10053 = n9936 ^ n9747;
  assign n10054 = n9937 & n10053;
  assign n10055 = n10054 ^ n9747;
  assign n10251 = n10250 ^ n10055;
  assign n10045 = n1404 & n6026;
  assign n10046 = x107 & n1514;
  assign n10047 = x108 & n1408;
  assign n10048 = ~n10046 & ~n10047;
  assign n10049 = x109 & n1517;
  assign n10050 = n10048 & ~n10049;
  assign n10051 = ~n10045 & n10050;
  assign n10052 = n10051 ^ x20;
  assign n10252 = n10251 ^ n10052;
  assign n10042 = n9938 ^ n9736;
  assign n10043 = ~n9939 & ~n10042;
  assign n10044 = n10043 ^ n9736;
  assign n10253 = n10252 ^ n10044;
  assign n10034 = n1098 & n6728;
  assign n10035 = x110 & n1198;
  assign n10036 = x111 & n1102;
  assign n10037 = ~n10035 & ~n10036;
  assign n10038 = x112 & n1201;
  assign n10039 = n10037 & ~n10038;
  assign n10040 = ~n10034 & n10039;
  assign n10041 = n10040 ^ x17;
  assign n10254 = n10253 ^ n10041;
  assign n10031 = n9940 ^ n9725;
  assign n10032 = n9941 & n10031;
  assign n10033 = n10032 ^ n9725;
  assign n10255 = n10254 ^ n10033;
  assign n10023 = n821 & n7481;
  assign n10024 = x113 & n898;
  assign n10025 = x115 & n901;
  assign n10026 = ~n10024 & ~n10025;
  assign n10027 = x114 & n824;
  assign n10028 = n10026 & ~n10027;
  assign n10029 = ~n10023 & n10028;
  assign n10030 = n10029 ^ x14;
  assign n10256 = n10255 ^ n10030;
  assign n10020 = n9942 ^ n9714;
  assign n10021 = ~n9943 & ~n10020;
  assign n10022 = n10021 ^ n9714;
  assign n10257 = n10256 ^ n10022;
  assign n10012 = n596 & n8265;
  assign n10013 = x116 & n673;
  assign n10014 = x118 & n676;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = x117 & n601;
  assign n10017 = n10015 & ~n10016;
  assign n10018 = ~n10012 & n10017;
  assign n10019 = n10018 ^ x11;
  assign n10258 = n10257 ^ n10019;
  assign n10009 = n9944 ^ n9703;
  assign n10010 = n9945 & n10009;
  assign n10011 = n10010 ^ n9703;
  assign n10259 = n10258 ^ n10011;
  assign n9999 = n9081 ^ x124;
  assign n10000 = n239 & n9999;
  assign n10001 = x122 & n249;
  assign n10002 = x123 & n242;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = x124 & n280;
  assign n10005 = n10003 & ~n10004;
  assign n10006 = ~n10000 & n10005;
  assign n10007 = n10006 ^ x5;
  assign n9991 = n399 & n9094;
  assign n9992 = x119 & n478;
  assign n9993 = x121 & n470;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = x120 & n402;
  assign n9996 = n9994 & ~n9995;
  assign n9997 = ~n9991 & n9996;
  assign n9998 = n9997 ^ x8;
  assign n10008 = n10007 ^ n9998;
  assign n10260 = n10259 ^ n10008;
  assign n9980 = x125 & ~x126;
  assign n9981 = ~n9673 & n9980;
  assign n9982 = ~x125 & x126;
  assign n9983 = ~n9675 & n9982;
  assign n9984 = ~n9981 & ~n9983;
  assign n9985 = n169 & n9984;
  assign n9986 = n9985 ^ x1;
  assign n9987 = n9986 ^ x127;
  assign n9972 = x126 ^ x2;
  assign n9973 = n9972 ^ x126;
  assign n9974 = n9972 ^ x125;
  assign n9975 = n9974 ^ n9972;
  assign n9976 = n9973 & ~n9975;
  assign n9977 = n9976 ^ n9972;
  assign n9978 = ~x1 & n9977;
  assign n9979 = n9978 ^ n9972;
  assign n9988 = n9987 ^ n9979;
  assign n9989 = ~x0 & n9988;
  assign n9990 = n9989 ^ n9987;
  assign n10261 = n10260 ^ n9990;
  assign n9969 = n9946 ^ n9699;
  assign n9970 = ~n9700 & n9969;
  assign n9971 = n9970 ^ n9946;
  assign n10262 = n10261 ^ n9971;
  assign n9966 = n9947 ^ n9659;
  assign n9967 = n9948 & ~n9966;
  assign n9968 = n9967 ^ n9659;
  assign n10263 = n10262 ^ n9968;
  assign n9963 = n9961 ^ n9949;
  assign n9964 = n9950 & n9963;
  assign n9965 = n9964 ^ n9961;
  assign n10264 = n10263 ^ n9965;
  assign n10518 = n956 & n7395;
  assign n10519 = x76 & n7400;
  assign n10520 = x75 & n7650;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = x77 & n7652;
  assign n10523 = n10521 & ~n10522;
  assign n10524 = ~n10518 & n10523;
  assign n10525 = n10524 ^ x53;
  assign n10515 = n10229 ^ n10166;
  assign n10516 = n10230 & n10515;
  assign n10517 = n10516 ^ n10166;
  assign n10526 = n10525 ^ n10517;
  assign n10507 = n10176 & n10185;
  assign n10508 = n10178 & ~n10186;
  assign n10509 = ~n10507 & ~n10508;
  assign n10497 = n321 & n9878;
  assign n10498 = x67 & n9881;
  assign n10499 = x66 & n9888;
  assign n10500 = ~n10498 & ~n10499;
  assign n10501 = n9296 & ~n9877;
  assign n10502 = x68 & n10501;
  assign n10503 = n10500 & ~n10502;
  assign n10504 = ~n10497 & n10503;
  assign n10505 = n10504 ^ x62;
  assign n10489 = x65 ^ x64;
  assign n10490 = n10489 ^ x65;
  assign n10491 = x65 ^ x63;
  assign n10492 = n10491 ^ x65;
  assign n10493 = n10490 & n10492;
  assign n10494 = n10493 ^ x65;
  assign n10495 = ~n10177 & n10494;
  assign n10496 = n10495 ^ x65;
  assign n10506 = n10505 ^ n10496;
  assign n10510 = n10509 ^ n10506;
  assign n10481 = n517 & n9002;
  assign n10482 = x69 & n9012;
  assign n10483 = x71 & n9557;
  assign n10484 = ~n10482 & ~n10483;
  assign n10485 = x70 & n9005;
  assign n10486 = n10484 & ~n10485;
  assign n10487 = ~n10481 & n10486;
  assign n10488 = n10487 ^ x59;
  assign n10511 = n10510 ^ n10488;
  assign n10478 = n10215 ^ n10195;
  assign n10479 = ~n10204 & n10478;
  assign n10480 = n10479 ^ n10215;
  assign n10512 = n10511 ^ n10480;
  assign n10470 = ~n721 & n8171;
  assign n10471 = x73 & n8174;
  assign n10472 = x72 & n8181;
  assign n10473 = ~n10471 & ~n10472;
  assign n10474 = x74 & n8732;
  assign n10475 = n10473 & ~n10474;
  assign n10476 = ~n10470 & n10475;
  assign n10477 = n10476 ^ x56;
  assign n10513 = n10512 ^ n10477;
  assign n10467 = n10227 ^ n10216;
  assign n10468 = ~n10228 & ~n10467;
  assign n10469 = n10468 ^ n10219;
  assign n10514 = n10513 ^ n10469;
  assign n10527 = n10526 ^ n10514;
  assign n10459 = n1242 & n6626;
  assign n10460 = x78 & n6884;
  assign n10461 = x79 & n6630;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = x80 & n6888;
  assign n10464 = n10462 & ~n10463;
  assign n10465 = ~n10459 & n10464;
  assign n10466 = n10465 ^ x50;
  assign n10528 = n10527 ^ n10466;
  assign n10456 = n10231 ^ n10159;
  assign n10457 = ~n10232 & ~n10456;
  assign n10458 = n10457 ^ n10163;
  assign n10529 = n10528 ^ n10458;
  assign n10448 = n1560 & n5942;
  assign n10449 = x81 & n6186;
  assign n10450 = x82 & n5947;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = x83 & n6406;
  assign n10453 = n10451 & ~n10452;
  assign n10454 = ~n10448 & n10453;
  assign n10455 = n10454 ^ x47;
  assign n10530 = n10529 ^ n10455;
  assign n10445 = n10233 ^ n10143;
  assign n10446 = n10234 & n10445;
  assign n10447 = n10446 ^ n10143;
  assign n10531 = n10530 ^ n10447;
  assign n10437 = n1920 & n5262;
  assign n10438 = x85 & n5266;
  assign n10439 = x86 & n5491;
  assign n10440 = ~n10438 & ~n10439;
  assign n10441 = x84 & n5488;
  assign n10442 = n10440 & ~n10441;
  assign n10443 = ~n10437 & n10442;
  assign n10444 = n10443 ^ x44;
  assign n10532 = n10531 ^ n10444;
  assign n10434 = n10235 ^ n10132;
  assign n10435 = ~n10236 & ~n10434;
  assign n10436 = n10435 ^ n10132;
  assign n10533 = n10532 ^ n10436;
  assign n10426 = n2310 & n4643;
  assign n10427 = x87 & n4653;
  assign n10428 = x88 & n4646;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = x89 & n5046;
  assign n10431 = n10429 & ~n10430;
  assign n10432 = ~n10426 & n10431;
  assign n10433 = n10432 ^ x41;
  assign n10534 = n10533 ^ n10433;
  assign n10423 = n10237 ^ n10121;
  assign n10424 = n10238 & n10423;
  assign n10425 = n10424 ^ n10121;
  assign n10535 = n10534 ^ n10425;
  assign n10415 = n2755 & n4040;
  assign n10416 = x90 & n4267;
  assign n10417 = x91 & n4044;
  assign n10418 = ~n10416 & ~n10417;
  assign n10419 = x92 & n4270;
  assign n10420 = n10418 & ~n10419;
  assign n10421 = ~n10415 & n10420;
  assign n10422 = n10421 ^ x38;
  assign n10536 = n10535 ^ n10422;
  assign n10412 = n10239 ^ n10110;
  assign n10413 = ~n10240 & ~n10412;
  assign n10414 = n10413 ^ n10110;
  assign n10537 = n10536 ^ n10414;
  assign n10404 = n3247 & n3522;
  assign n10405 = x93 & n3699;
  assign n10406 = x94 & n3526;
  assign n10407 = ~n10405 & ~n10406;
  assign n10408 = x95 & n3701;
  assign n10409 = n10407 & ~n10408;
  assign n10410 = ~n10404 & n10409;
  assign n10411 = n10410 ^ x35;
  assign n10538 = n10537 ^ n10411;
  assign n10401 = n10241 ^ n10099;
  assign n10402 = n10242 & n10401;
  assign n10403 = n10402 ^ n10099;
  assign n10539 = n10538 ^ n10403;
  assign n10393 = n3009 & n3763;
  assign n10394 = x96 & n3181;
  assign n10395 = x97 & n3013;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = x98 & n3183;
  assign n10398 = n10396 & ~n10397;
  assign n10399 = ~n10393 & n10398;
  assign n10400 = n10399 ^ x32;
  assign n10540 = n10539 ^ n10400;
  assign n10390 = n10243 ^ n10088;
  assign n10391 = ~n10244 & ~n10390;
  assign n10392 = n10391 ^ n10088;
  assign n10541 = n10540 ^ n10392;
  assign n10382 = n2527 & n4323;
  assign n10383 = x100 & n2530;
  assign n10384 = x99 & n2690;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = x101 & n2693;
  assign n10387 = n10385 & ~n10386;
  assign n10388 = ~n10382 & n10387;
  assign n10389 = n10388 ^ x29;
  assign n10542 = n10541 ^ n10389;
  assign n10379 = n10245 ^ n10077;
  assign n10380 = n10246 & n10379;
  assign n10381 = n10380 ^ n10077;
  assign n10543 = n10542 ^ n10381;
  assign n10371 = n2102 & n4912;
  assign n10372 = x102 & n2112;
  assign n10373 = x103 & n2105;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = x104 & n2381;
  assign n10376 = n10374 & ~n10375;
  assign n10377 = ~n10371 & n10376;
  assign n10378 = n10377 ^ x26;
  assign n10544 = n10543 ^ n10378;
  assign n10368 = n10247 ^ n10066;
  assign n10369 = ~n10248 & ~n10368;
  assign n10370 = n10369 ^ n10066;
  assign n10545 = n10544 ^ n10370;
  assign n10360 = n1746 & n5578;
  assign n10361 = x106 & n1750;
  assign n10362 = x105 & n1871;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = x107 & n1873;
  assign n10365 = n10363 & ~n10364;
  assign n10366 = ~n10360 & n10365;
  assign n10367 = n10366 ^ x23;
  assign n10546 = n10545 ^ n10367;
  assign n10357 = n10249 ^ n10055;
  assign n10358 = n10250 & n10357;
  assign n10359 = n10358 ^ n10055;
  assign n10547 = n10546 ^ n10359;
  assign n10349 = n1404 & n6250;
  assign n10350 = x109 & n1408;
  assign n10351 = x108 & n1514;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = x110 & n1517;
  assign n10354 = n10352 & ~n10353;
  assign n10355 = ~n10349 & n10354;
  assign n10356 = n10355 ^ x20;
  assign n10548 = n10547 ^ n10356;
  assign n10346 = n10251 ^ n10044;
  assign n10347 = ~n10252 & ~n10346;
  assign n10348 = n10347 ^ n10044;
  assign n10549 = n10548 ^ n10348;
  assign n10338 = n1098 & n6975;
  assign n10339 = x111 & n1198;
  assign n10340 = x112 & n1102;
  assign n10341 = ~n10339 & ~n10340;
  assign n10342 = x113 & n1201;
  assign n10343 = n10341 & ~n10342;
  assign n10344 = ~n10338 & n10343;
  assign n10345 = n10344 ^ x17;
  assign n10550 = n10549 ^ n10345;
  assign n10335 = n10253 ^ n10033;
  assign n10336 = n10254 & n10335;
  assign n10337 = n10336 ^ n10033;
  assign n10551 = n10550 ^ n10337;
  assign n10327 = n821 & n7730;
  assign n10328 = x115 & n824;
  assign n10329 = x114 & n898;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = x116 & n901;
  assign n10332 = n10330 & ~n10331;
  assign n10333 = ~n10327 & n10332;
  assign n10334 = n10333 ^ x14;
  assign n10552 = n10551 ^ n10334;
  assign n10324 = n10255 ^ n10022;
  assign n10325 = ~n10256 & ~n10324;
  assign n10326 = n10325 ^ n10022;
  assign n10553 = n10552 ^ n10326;
  assign n10316 = n596 & n8542;
  assign n10317 = x117 & n673;
  assign n10318 = x118 & n601;
  assign n10319 = ~n10317 & ~n10318;
  assign n10320 = x119 & n676;
  assign n10321 = n10319 & ~n10320;
  assign n10322 = ~n10316 & n10321;
  assign n10323 = n10322 ^ x11;
  assign n10554 = n10553 ^ n10323;
  assign n10313 = n10257 ^ n10011;
  assign n10314 = n10258 & n10313;
  assign n10315 = n10314 ^ n10011;
  assign n10555 = n10554 ^ n10315;
  assign n10302 = x125 ^ x124;
  assign n10303 = n10302 ^ n9365;
  assign n10304 = n239 & n10303;
  assign n10305 = x123 & n249;
  assign n10306 = x125 & n280;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = x124 & n242;
  assign n10309 = n10307 & ~n10308;
  assign n10310 = ~n10304 & n10309;
  assign n10311 = n10310 ^ x5;
  assign n10294 = n399 & n9387;
  assign n10295 = x120 & n478;
  assign n10296 = x121 & n402;
  assign n10297 = ~n10295 & ~n10296;
  assign n10298 = x122 & n470;
  assign n10299 = n10297 & ~n10298;
  assign n10300 = ~n10294 & n10299;
  assign n10301 = n10300 ^ x8;
  assign n10312 = n10311 ^ n10301;
  assign n10556 = n10555 ^ n10312;
  assign n10274 = ~x1 & x126;
  assign n10275 = x2 & ~x127;
  assign n10276 = ~n10274 & n10275;
  assign n10277 = ~x126 & x127;
  assign n10278 = ~n9981 & n10277;
  assign n10279 = x126 & ~x127;
  assign n10280 = ~n9983 & n10279;
  assign n10281 = ~n10278 & ~n10280;
  assign n10282 = n169 & n10281;
  assign n10283 = n10282 ^ x1;
  assign n10284 = n10283 ^ x0;
  assign n10285 = n10284 ^ n10283;
  assign n10286 = x127 ^ x126;
  assign n10287 = ~n9973 & ~n10286;
  assign n10288 = n10287 ^ x126;
  assign n10289 = n169 & ~n10288;
  assign n10290 = n10289 ^ n10283;
  assign n10291 = ~n10285 & n10290;
  assign n10292 = n10291 ^ n10283;
  assign n10293 = ~n10276 & ~n10292;
  assign n10557 = n10556 ^ n10293;
  assign n10271 = n10259 ^ n10007;
  assign n10272 = ~n10008 & n10271;
  assign n10273 = n10272 ^ n10259;
  assign n10558 = n10557 ^ n10273;
  assign n10268 = n9990 ^ n9971;
  assign n10269 = ~n10261 & n10268;
  assign n10270 = n10269 ^ n10260;
  assign n10559 = n10558 ^ n10270;
  assign n10265 = n9968 ^ n9965;
  assign n10266 = ~n10263 & ~n10265;
  assign n10267 = n10266 ^ n9965;
  assign n10560 = n10559 ^ n10267;
  assign n10842 = n10555 ^ n10311;
  assign n10843 = ~n10312 & ~n10842;
  assign n10844 = n10843 ^ n10555;
  assign n10828 = n169 ^ x127;
  assign n10829 = x2 ^ x0;
  assign n10830 = n10829 ^ x2;
  assign n10831 = n10278 ^ x2;
  assign n10832 = n10830 & ~n10831;
  assign n10833 = n10832 ^ x2;
  assign n10834 = n10833 ^ n169;
  assign n10835 = n10828 & n10834;
  assign n10836 = n10835 ^ n10832;
  assign n10837 = n10836 ^ x2;
  assign n10838 = n10837 ^ x127;
  assign n10839 = n169 & n10838;
  assign n10840 = n10839 ^ n169;
  assign n10841 = n10840 ^ x2;
  assign n10845 = n10844 ^ n10841;
  assign n10789 = n1041 & n7395;
  assign n10790 = x77 & n7400;
  assign n10791 = x76 & n7650;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = x78 & n7652;
  assign n10794 = n10792 & ~n10793;
  assign n10795 = ~n10789 & n10794;
  assign n10796 = n10795 ^ x53;
  assign n10786 = n10525 ^ n10514;
  assign n10787 = ~n10526 & ~n10786;
  assign n10788 = n10787 ^ n10517;
  assign n10797 = n10796 ^ n10788;
  assign n10776 = n789 & n8171;
  assign n10777 = x74 & n8174;
  assign n10778 = x73 & n8181;
  assign n10779 = ~n10777 & ~n10778;
  assign n10780 = x75 & n8732;
  assign n10781 = n10779 & ~n10780;
  assign n10782 = ~n10776 & n10781;
  assign n10783 = n10782 ^ x56;
  assign n10773 = n10512 ^ n10469;
  assign n10774 = n10513 & n10773;
  assign n10775 = n10774 ^ n10469;
  assign n10784 = n10783 ^ n10775;
  assign n10761 = x66 ^ x65;
  assign n10762 = n10761 ^ x66;
  assign n10763 = x66 ^ x63;
  assign n10764 = n10763 ^ x66;
  assign n10765 = n10762 & n10764;
  assign n10766 = n10765 ^ x66;
  assign n10767 = ~n10177 & n10766;
  assign n10768 = n10767 ^ x66;
  assign n10758 = n10509 ^ n10505;
  assign n10759 = n10506 & n10758;
  assign n10760 = n10759 ^ n10509;
  assign n10769 = n10768 ^ n10760;
  assign n10750 = n420 & n9878;
  assign n10751 = x68 & n9881;
  assign n10752 = x67 & n9888;
  assign n10753 = ~n10751 & ~n10752;
  assign n10754 = x69 & n10501;
  assign n10755 = n10753 & ~n10754;
  assign n10756 = ~n10750 & n10755;
  assign n10757 = n10756 ^ x62;
  assign n10770 = n10769 ^ n10757;
  assign n10742 = n575 & n9002;
  assign n10743 = x70 & n9012;
  assign n10744 = x71 & n9005;
  assign n10745 = ~n10743 & ~n10744;
  assign n10746 = x72 & n9557;
  assign n10747 = n10745 & ~n10746;
  assign n10748 = ~n10742 & n10747;
  assign n10749 = n10748 ^ x59;
  assign n10771 = n10770 ^ n10749;
  assign n10739 = n10510 ^ n10480;
  assign n10740 = n10511 & ~n10739;
  assign n10741 = n10740 ^ n10480;
  assign n10772 = n10771 ^ n10741;
  assign n10785 = n10784 ^ n10772;
  assign n10798 = n10797 ^ n10785;
  assign n10731 = n1340 & n6626;
  assign n10732 = x79 & n6884;
  assign n10733 = x80 & n6630;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = x81 & n6888;
  assign n10736 = n10734 & ~n10735;
  assign n10737 = ~n10731 & n10736;
  assign n10738 = n10737 ^ x50;
  assign n10799 = n10798 ^ n10738;
  assign n10728 = n10527 ^ n10458;
  assign n10729 = n10528 & n10728;
  assign n10730 = n10729 ^ n10458;
  assign n10800 = n10799 ^ n10730;
  assign n10720 = n1667 & n5942;
  assign n10721 = x82 & n6186;
  assign n10722 = x84 & n6406;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = x83 & n5947;
  assign n10725 = n10723 & ~n10724;
  assign n10726 = ~n10720 & n10725;
  assign n10727 = n10726 ^ x47;
  assign n10801 = n10800 ^ n10727;
  assign n10717 = n10529 ^ n10447;
  assign n10718 = ~n10530 & ~n10717;
  assign n10719 = n10718 ^ n10447;
  assign n10802 = n10801 ^ n10719;
  assign n10709 = n2039 & n5262;
  assign n10710 = x85 & n5488;
  assign n10711 = x86 & n5266;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = x87 & n5491;
  assign n10714 = n10712 & ~n10713;
  assign n10715 = ~n10709 & n10714;
  assign n10716 = n10715 ^ x44;
  assign n10803 = n10802 ^ n10716;
  assign n10706 = n10531 ^ n10436;
  assign n10707 = n10532 & n10706;
  assign n10708 = n10707 ^ n10436;
  assign n10804 = n10803 ^ n10708;
  assign n10698 = n2448 & n4643;
  assign n10699 = x88 & n4653;
  assign n10700 = x90 & n5046;
  assign n10701 = ~n10699 & ~n10700;
  assign n10702 = x89 & n4646;
  assign n10703 = n10701 & ~n10702;
  assign n10704 = ~n10698 & n10703;
  assign n10705 = n10704 ^ x41;
  assign n10805 = n10804 ^ n10705;
  assign n10695 = n10533 ^ n10425;
  assign n10696 = ~n10534 & ~n10695;
  assign n10697 = n10696 ^ n10425;
  assign n10806 = n10805 ^ n10697;
  assign n10687 = n2901 & n4040;
  assign n10688 = x91 & n4267;
  assign n10689 = x93 & n4270;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = x92 & n4044;
  assign n10692 = n10690 & ~n10691;
  assign n10693 = ~n10687 & n10692;
  assign n10694 = n10693 ^ x38;
  assign n10807 = n10806 ^ n10694;
  assign n10684 = n10535 ^ n10414;
  assign n10685 = n10536 & n10684;
  assign n10686 = n10685 ^ n10414;
  assign n10808 = n10807 ^ n10686;
  assign n10676 = n3403 & n3522;
  assign n10677 = x94 & n3699;
  assign n10678 = x96 & n3701;
  assign n10679 = ~n10677 & ~n10678;
  assign n10680 = x95 & n3526;
  assign n10681 = n10679 & ~n10680;
  assign n10682 = ~n10676 & n10681;
  assign n10683 = n10682 ^ x35;
  assign n10809 = n10808 ^ n10683;
  assign n10673 = n10537 ^ n10403;
  assign n10674 = ~n10538 & ~n10673;
  assign n10675 = n10674 ^ n10403;
  assign n10810 = n10809 ^ n10675;
  assign n10665 = n3009 & n3943;
  assign n10666 = x97 & n3181;
  assign n10667 = x98 & n3013;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = x99 & n3183;
  assign n10670 = n10668 & ~n10669;
  assign n10671 = ~n10665 & n10670;
  assign n10672 = n10671 ^ x32;
  assign n10811 = n10810 ^ n10672;
  assign n10662 = n10539 ^ n10392;
  assign n10663 = n10540 & n10662;
  assign n10664 = n10663 ^ n10392;
  assign n10812 = n10811 ^ n10664;
  assign n10654 = n2527 & n4509;
  assign n10655 = x101 & n2530;
  assign n10656 = x100 & n2690;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = x102 & n2693;
  assign n10659 = n10657 & ~n10658;
  assign n10660 = ~n10654 & n10659;
  assign n10661 = n10660 ^ x29;
  assign n10813 = n10812 ^ n10661;
  assign n10651 = n10541 ^ n10381;
  assign n10652 = ~n10542 & ~n10651;
  assign n10653 = n10652 ^ n10381;
  assign n10814 = n10813 ^ n10653;
  assign n10643 = n2102 & n5117;
  assign n10644 = x103 & n2112;
  assign n10645 = x105 & n2381;
  assign n10646 = ~n10644 & ~n10645;
  assign n10647 = x104 & n2105;
  assign n10648 = n10646 & ~n10647;
  assign n10649 = ~n10643 & n10648;
  assign n10650 = n10649 ^ x26;
  assign n10815 = n10814 ^ n10650;
  assign n10640 = n10543 ^ n10370;
  assign n10641 = n10544 & n10640;
  assign n10642 = n10641 ^ n10370;
  assign n10816 = n10815 ^ n10642;
  assign n10632 = n1746 & n5792;
  assign n10633 = x106 & n1871;
  assign n10634 = x108 & n1873;
  assign n10635 = ~n10633 & ~n10634;
  assign n10636 = x107 & n1750;
  assign n10637 = n10635 & ~n10636;
  assign n10638 = ~n10632 & n10637;
  assign n10639 = n10638 ^ x23;
  assign n10817 = n10816 ^ n10639;
  assign n10629 = n10545 ^ n10359;
  assign n10630 = ~n10546 & ~n10629;
  assign n10631 = n10630 ^ n10359;
  assign n10818 = n10817 ^ n10631;
  assign n10621 = n1404 & n6478;
  assign n10622 = x109 & n1514;
  assign n10623 = x110 & n1408;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 = x111 & n1517;
  assign n10626 = n10624 & ~n10625;
  assign n10627 = ~n10621 & n10626;
  assign n10628 = n10627 ^ x20;
  assign n10819 = n10818 ^ n10628;
  assign n10618 = n10547 ^ n10348;
  assign n10619 = n10548 & n10618;
  assign n10620 = n10619 ^ n10348;
  assign n10820 = n10819 ^ n10620;
  assign n10610 = n1098 & n7220;
  assign n10611 = x113 & n1102;
  assign n10612 = x112 & n1198;
  assign n10613 = ~n10611 & ~n10612;
  assign n10614 = x114 & n1201;
  assign n10615 = n10613 & ~n10614;
  assign n10616 = ~n10610 & n10615;
  assign n10617 = n10616 ^ x17;
  assign n10821 = n10820 ^ n10617;
  assign n10607 = n10549 ^ n10337;
  assign n10608 = ~n10550 & ~n10607;
  assign n10609 = n10608 ^ n10337;
  assign n10822 = n10821 ^ n10609;
  assign n10599 = n821 & n7987;
  assign n10600 = x115 & n898;
  assign n10601 = x116 & n824;
  assign n10602 = ~n10600 & ~n10601;
  assign n10603 = x117 & n901;
  assign n10604 = n10602 & ~n10603;
  assign n10605 = ~n10599 & n10604;
  assign n10606 = n10605 ^ x14;
  assign n10823 = n10822 ^ n10606;
  assign n10596 = n10551 ^ n10326;
  assign n10597 = n10552 & n10596;
  assign n10598 = n10597 ^ n10326;
  assign n10824 = n10823 ^ n10598;
  assign n10587 = n399 & n9691;
  assign n10588 = x121 & n478;
  assign n10589 = x123 & n470;
  assign n10590 = ~n10588 & ~n10589;
  assign n10591 = x122 & n402;
  assign n10592 = n10590 & ~n10591;
  assign n10593 = ~n10587 & n10592;
  assign n10594 = n10593 ^ x8;
  assign n10579 = n596 & n8820;
  assign n10580 = x119 & n601;
  assign n10581 = x118 & n673;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = x120 & n676;
  assign n10584 = n10582 & ~n10583;
  assign n10585 = ~n10579 & n10584;
  assign n10586 = n10585 ^ x11;
  assign n10595 = n10594 ^ n10586;
  assign n10825 = n10824 ^ n10595;
  assign n10570 = n9676 ^ x126;
  assign n10571 = n239 & ~n10570;
  assign n10572 = x124 & n249;
  assign n10573 = x125 & n242;
  assign n10574 = ~n10572 & ~n10573;
  assign n10575 = x126 & n280;
  assign n10576 = n10574 & ~n10575;
  assign n10577 = ~n10571 & n10576;
  assign n10578 = n10577 ^ x5;
  assign n10826 = n10825 ^ n10578;
  assign n10567 = n10553 ^ n10315;
  assign n10568 = ~n10554 & ~n10567;
  assign n10569 = n10568 ^ n10315;
  assign n10827 = n10826 ^ n10569;
  assign n10846 = n10845 ^ n10827;
  assign n10564 = n10293 ^ n10273;
  assign n10565 = ~n10557 & ~n10564;
  assign n10566 = n10565 ^ n10556;
  assign n10847 = n10846 ^ n10566;
  assign n10561 = n10558 ^ n10267;
  assign n10562 = n10559 & ~n10561;
  assign n10563 = n10562 ^ n10267;
  assign n10848 = n10847 ^ n10563;
  assign n11073 = ~n653 & n9002;
  assign n11074 = x72 & n9005;
  assign n11075 = x71 & n9012;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = x73 & n9557;
  assign n11078 = n11076 & ~n11077;
  assign n11079 = ~n11073 & n11078;
  assign n11080 = n11079 ^ x59;
  assign n11065 = n458 & n9878;
  assign n11066 = x68 & n9888;
  assign n11067 = x70 & n10501;
  assign n11068 = ~n11066 & ~n11067;
  assign n11069 = x69 & n9881;
  assign n11070 = n11068 & ~n11069;
  assign n11071 = ~n11065 & n11070;
  assign n11060 = x63 & x67;
  assign n11057 = x67 ^ x66;
  assign n11058 = ~x63 & n11057;
  assign n11059 = n11058 ^ x66;
  assign n11061 = n11060 ^ n11059;
  assign n11062 = ~x62 & ~n11061;
  assign n11063 = n11062 ^ n11059;
  assign n11064 = n11063 ^ x2;
  assign n11072 = n11071 ^ n11064;
  assign n11081 = n11080 ^ n11072;
  assign n11054 = n10768 ^ n10757;
  assign n11055 = ~n10769 & n11054;
  assign n11056 = n11055 ^ n10760;
  assign n11082 = n11081 ^ n11056;
  assign n11046 = n870 & n8171;
  assign n11047 = x74 & n8181;
  assign n11048 = x75 & n8174;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = x76 & n8732;
  assign n11051 = n11049 & ~n11050;
  assign n11052 = ~n11046 & n11051;
  assign n11053 = n11052 ^ x56;
  assign n11083 = n11082 ^ n11053;
  assign n11043 = n10770 ^ n10741;
  assign n11044 = n10771 & ~n11043;
  assign n11045 = n11044 ^ n10741;
  assign n11084 = n11083 ^ n11045;
  assign n11035 = n1149 & n7395;
  assign n11036 = x78 & n7400;
  assign n11037 = x77 & n7650;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = x79 & n7652;
  assign n11040 = n11038 & ~n11039;
  assign n11041 = ~n11035 & n11040;
  assign n11042 = n11041 ^ x53;
  assign n11085 = n11084 ^ n11042;
  assign n11032 = n10783 ^ n10772;
  assign n11033 = ~n10784 & n11032;
  assign n11034 = n11033 ^ n10775;
  assign n11086 = n11085 ^ n11034;
  assign n11024 = n1454 & n6626;
  assign n11025 = x80 & n6884;
  assign n11026 = x81 & n6630;
  assign n11027 = ~n11025 & ~n11026;
  assign n11028 = x82 & n6888;
  assign n11029 = n11027 & ~n11028;
  assign n11030 = ~n11024 & n11029;
  assign n11031 = n11030 ^ x50;
  assign n11087 = n11086 ^ n11031;
  assign n11021 = n10796 ^ n10785;
  assign n11022 = ~n10797 & ~n11021;
  assign n11023 = n11022 ^ n10788;
  assign n11088 = n11087 ^ n11023;
  assign n11013 = n1801 & n5942;
  assign n11014 = x83 & n6186;
  assign n11015 = x85 & n6406;
  assign n11016 = ~n11014 & ~n11015;
  assign n11017 = x84 & n5947;
  assign n11018 = n11016 & ~n11017;
  assign n11019 = ~n11013 & n11018;
  assign n11020 = n11019 ^ x47;
  assign n11089 = n11088 ^ n11020;
  assign n11010 = n10798 ^ n10730;
  assign n11011 = n10799 & n11010;
  assign n11012 = n11011 ^ n10730;
  assign n11090 = n11089 ^ n11012;
  assign n11002 = n2176 & n5262;
  assign n11003 = x86 & n5488;
  assign n11004 = x88 & n5491;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = x87 & n5266;
  assign n11007 = n11005 & ~n11006;
  assign n11008 = ~n11002 & n11007;
  assign n11009 = n11008 ^ x44;
  assign n11091 = n11090 ^ n11009;
  assign n10999 = n10800 ^ n10719;
  assign n11000 = ~n10801 & ~n10999;
  assign n11001 = n11000 ^ n10719;
  assign n11092 = n11091 ^ n11001;
  assign n10991 = n2607 & n4643;
  assign n10992 = x89 & n4653;
  assign n10993 = x90 & n4646;
  assign n10994 = ~n10992 & ~n10993;
  assign n10995 = x91 & n5046;
  assign n10996 = n10994 & ~n10995;
  assign n10997 = ~n10991 & n10996;
  assign n10998 = n10997 ^ x41;
  assign n11093 = n11092 ^ n10998;
  assign n10988 = n10802 ^ n10708;
  assign n10989 = n10803 & n10988;
  assign n10990 = n10989 ^ n10708;
  assign n11094 = n11093 ^ n10990;
  assign n10980 = n3078 & n4040;
  assign n10981 = x93 & n4044;
  assign n10982 = x92 & n4267;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = x94 & n4270;
  assign n10985 = n10983 & ~n10984;
  assign n10986 = ~n10980 & n10985;
  assign n10987 = n10986 ^ x38;
  assign n11095 = n11094 ^ n10987;
  assign n10977 = n10804 ^ n10697;
  assign n10978 = ~n10805 & ~n10977;
  assign n10979 = n10978 ^ n10697;
  assign n11096 = n11095 ^ n10979;
  assign n10969 = n3522 & n3585;
  assign n10970 = x95 & n3699;
  assign n10971 = x96 & n3526;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = x97 & n3701;
  assign n10974 = n10972 & ~n10973;
  assign n10975 = ~n10969 & n10974;
  assign n10976 = n10975 ^ x35;
  assign n11097 = n11096 ^ n10976;
  assign n10966 = n10806 ^ n10686;
  assign n10967 = n10807 & n10966;
  assign n10968 = n10967 ^ n10686;
  assign n11098 = n11097 ^ n10968;
  assign n10958 = n3009 & n4141;
  assign n10959 = x99 & n3013;
  assign n10960 = x98 & n3181;
  assign n10961 = ~n10959 & ~n10960;
  assign n10962 = x100 & n3183;
  assign n10963 = n10961 & ~n10962;
  assign n10964 = ~n10958 & n10963;
  assign n10965 = n10964 ^ x32;
  assign n11099 = n11098 ^ n10965;
  assign n10955 = n10808 ^ n10675;
  assign n10956 = ~n10809 & ~n10955;
  assign n10957 = n10956 ^ n10675;
  assign n11100 = n11099 ^ n10957;
  assign n10947 = n2527 & n4718;
  assign n10948 = x101 & n2690;
  assign n10949 = x103 & n2693;
  assign n10950 = ~n10948 & ~n10949;
  assign n10951 = x102 & n2530;
  assign n10952 = n10950 & ~n10951;
  assign n10953 = ~n10947 & n10952;
  assign n10954 = n10953 ^ x29;
  assign n11101 = n11100 ^ n10954;
  assign n10944 = n10810 ^ n10664;
  assign n10945 = n10811 & n10944;
  assign n10946 = n10945 ^ n10664;
  assign n11102 = n11101 ^ n10946;
  assign n10936 = n2102 & n5351;
  assign n10937 = x104 & n2112;
  assign n10938 = x106 & n2381;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = x105 & n2105;
  assign n10941 = n10939 & ~n10940;
  assign n10942 = ~n10936 & n10941;
  assign n10943 = n10942 ^ x26;
  assign n11103 = n11102 ^ n10943;
  assign n10933 = n10812 ^ n10653;
  assign n10934 = ~n10813 & ~n10933;
  assign n10935 = n10934 ^ n10653;
  assign n11104 = n11103 ^ n10935;
  assign n10925 = n1746 & n6026;
  assign n10926 = x107 & n1871;
  assign n10927 = x108 & n1750;
  assign n10928 = ~n10926 & ~n10927;
  assign n10929 = x109 & n1873;
  assign n10930 = n10928 & ~n10929;
  assign n10931 = ~n10925 & n10930;
  assign n10932 = n10931 ^ x23;
  assign n11105 = n11104 ^ n10932;
  assign n10922 = n10814 ^ n10642;
  assign n10923 = n10815 & n10922;
  assign n10924 = n10923 ^ n10642;
  assign n11106 = n11105 ^ n10924;
  assign n10914 = n1404 & n6728;
  assign n10915 = x110 & n1514;
  assign n10916 = x111 & n1408;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = x112 & n1517;
  assign n10919 = n10917 & ~n10918;
  assign n10920 = ~n10914 & n10919;
  assign n10921 = n10920 ^ x20;
  assign n11107 = n11106 ^ n10921;
  assign n10911 = n10816 ^ n10631;
  assign n10912 = ~n10817 & ~n10911;
  assign n10913 = n10912 ^ n10631;
  assign n11108 = n11107 ^ n10913;
  assign n10903 = n1098 & n7481;
  assign n10904 = x114 & n1102;
  assign n10905 = x113 & n1198;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = x115 & n1201;
  assign n10908 = n10906 & ~n10907;
  assign n10909 = ~n10903 & n10908;
  assign n10910 = n10909 ^ x17;
  assign n11109 = n11108 ^ n10910;
  assign n10900 = n10818 ^ n10620;
  assign n10901 = n10819 & n10900;
  assign n10902 = n10901 ^ n10620;
  assign n11110 = n11109 ^ n10902;
  assign n10892 = n821 & n8265;
  assign n10893 = x116 & n898;
  assign n10894 = x117 & n824;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = x118 & n901;
  assign n10897 = n10895 & ~n10896;
  assign n10898 = ~n10892 & n10897;
  assign n10899 = n10898 ^ x14;
  assign n11111 = n11110 ^ n10899;
  assign n10889 = n10820 ^ n10609;
  assign n10890 = ~n10821 & ~n10889;
  assign n10891 = n10890 ^ n10609;
  assign n11112 = n11111 ^ n10891;
  assign n10881 = n596 & n9094;
  assign n10882 = x119 & n673;
  assign n10883 = x121 & n676;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = x120 & n601;
  assign n10886 = n10884 & ~n10885;
  assign n10887 = ~n10881 & n10886;
  assign n10888 = n10887 ^ x11;
  assign n11113 = n11112 ^ n10888;
  assign n10878 = n10822 ^ n10598;
  assign n10879 = n10823 & n10878;
  assign n10880 = n10879 ^ n10598;
  assign n11114 = n11113 ^ n10880;
  assign n10875 = n10824 ^ n10594;
  assign n10876 = ~n10595 & n10875;
  assign n10877 = n10876 ^ n10824;
  assign n11115 = n11114 ^ n10877;
  assign n10867 = n399 & n9999;
  assign n10868 = x122 & n478;
  assign n10869 = x124 & n470;
  assign n10870 = ~n10868 & ~n10869;
  assign n10871 = x123 & n402;
  assign n10872 = n10870 & ~n10871;
  assign n10873 = ~n10867 & n10872;
  assign n10874 = n10873 ^ x8;
  assign n11116 = n11115 ^ n10874;
  assign n10864 = n10825 ^ n10569;
  assign n10865 = ~n10826 & ~n10864;
  assign n10866 = n10865 ^ n10569;
  assign n11117 = n11116 ^ n10866;
  assign n10855 = n9984 ^ x127;
  assign n10856 = n239 & ~n10855;
  assign n10857 = x125 & n249;
  assign n10858 = x127 & n280;
  assign n10859 = ~n10857 & ~n10858;
  assign n10860 = x126 & n242;
  assign n10861 = n10859 & ~n10860;
  assign n10862 = ~n10856 & n10861;
  assign n10863 = n10862 ^ x5;
  assign n11118 = n11117 ^ n10863;
  assign n10852 = n10841 ^ n10827;
  assign n10853 = n10845 & ~n10852;
  assign n10854 = n10853 ^ n10844;
  assign n11119 = n11118 ^ n10854;
  assign n10849 = n10846 ^ n10563;
  assign n10850 = ~n10847 & ~n10849;
  assign n10851 = n10850 ^ n10563;
  assign n11120 = n11119 ^ n10851;
  assign n11355 = n1560 & n6626;
  assign n11356 = x81 & n6884;
  assign n11357 = x83 & n6888;
  assign n11358 = ~n11356 & ~n11357;
  assign n11359 = x82 & n6630;
  assign n11360 = n11358 & ~n11359;
  assign n11361 = ~n11355 & n11360;
  assign n11362 = n11361 ^ x50;
  assign n11352 = n11084 ^ n11034;
  assign n11353 = n11085 & n11352;
  assign n11354 = n11353 ^ n11034;
  assign n11363 = n11362 ^ n11354;
  assign n11342 = n1242 & n7395;
  assign n11343 = x79 & n7400;
  assign n11344 = x80 & n7652;
  assign n11345 = ~n11343 & ~n11344;
  assign n11346 = x78 & n7650;
  assign n11347 = n11345 & ~n11346;
  assign n11348 = ~n11342 & n11347;
  assign n11349 = n11348 ^ x53;
  assign n11332 = n956 & n8171;
  assign n11333 = x75 & n8181;
  assign n11334 = x77 & n8732;
  assign n11335 = ~n11333 & ~n11334;
  assign n11336 = x76 & n8174;
  assign n11337 = n11335 & ~n11336;
  assign n11338 = ~n11332 & n11337;
  assign n11339 = n11338 ^ x56;
  assign n11322 = n517 & n9878;
  assign n11323 = x69 & n9888;
  assign n11324 = x71 & n10501;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = x70 & n9881;
  assign n11327 = n11325 & ~n11326;
  assign n11328 = ~n11322 & n11327;
  assign n11317 = x63 & x68;
  assign n11314 = x68 ^ x67;
  assign n11315 = ~x63 & n11314;
  assign n11316 = n11315 ^ x67;
  assign n11318 = n11317 ^ n11316;
  assign n11319 = ~x62 & ~n11318;
  assign n11320 = n11319 ^ n11316;
  assign n11321 = n11320 ^ x2;
  assign n11329 = n11328 ^ n11321;
  assign n11304 = n11071 ^ x2;
  assign n11308 = n11059 ^ x2;
  assign n11309 = n11304 & n11308;
  assign n11310 = n11309 ^ x2;
  assign n11305 = n11060 ^ x2;
  assign n11306 = ~n11304 & n11305;
  assign n11307 = n11306 ^ x2;
  assign n11311 = n11310 ^ n11307;
  assign n11312 = ~x62 & n11311;
  assign n11313 = n11312 ^ n11310;
  assign n11330 = n11329 ^ n11313;
  assign n11296 = ~n721 & n9002;
  assign n11297 = x73 & n9005;
  assign n11298 = x72 & n9012;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = x74 & n9557;
  assign n11301 = n11299 & ~n11300;
  assign n11302 = ~n11296 & n11301;
  assign n11303 = n11302 ^ x59;
  assign n11331 = n11330 ^ n11303;
  assign n11340 = n11339 ^ n11331;
  assign n11293 = n11080 ^ n11056;
  assign n11294 = n11081 & n11293;
  assign n11295 = n11294 ^ n11056;
  assign n11341 = n11340 ^ n11295;
  assign n11350 = n11349 ^ n11341;
  assign n11290 = n11082 ^ n11045;
  assign n11291 = n11083 & ~n11290;
  assign n11292 = n11291 ^ n11045;
  assign n11351 = n11350 ^ n11292;
  assign n11364 = n11363 ^ n11351;
  assign n11282 = n1920 & n5942;
  assign n11283 = x84 & n6186;
  assign n11284 = x86 & n6406;
  assign n11285 = ~n11283 & ~n11284;
  assign n11286 = x85 & n5947;
  assign n11287 = n11285 & ~n11286;
  assign n11288 = ~n11282 & n11287;
  assign n11289 = n11288 ^ x47;
  assign n11365 = n11364 ^ n11289;
  assign n11279 = n11086 ^ n11023;
  assign n11280 = ~n11087 & ~n11279;
  assign n11281 = n11280 ^ n11023;
  assign n11366 = n11365 ^ n11281;
  assign n11271 = n2310 & n5262;
  assign n11272 = x87 & n5488;
  assign n11273 = x88 & n5266;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = x89 & n5491;
  assign n11276 = n11274 & ~n11275;
  assign n11277 = ~n11271 & n11276;
  assign n11278 = n11277 ^ x44;
  assign n11367 = n11366 ^ n11278;
  assign n11268 = n11088 ^ n11012;
  assign n11269 = n11089 & n11268;
  assign n11270 = n11269 ^ n11012;
  assign n11368 = n11367 ^ n11270;
  assign n11260 = n2755 & n4643;
  assign n11261 = x90 & n4653;
  assign n11262 = x91 & n4646;
  assign n11263 = ~n11261 & ~n11262;
  assign n11264 = x92 & n5046;
  assign n11265 = n11263 & ~n11264;
  assign n11266 = ~n11260 & n11265;
  assign n11267 = n11266 ^ x41;
  assign n11369 = n11368 ^ n11267;
  assign n11257 = n11090 ^ n11001;
  assign n11258 = ~n11091 & ~n11257;
  assign n11259 = n11258 ^ n11001;
  assign n11370 = n11369 ^ n11259;
  assign n11249 = n3247 & n4040;
  assign n11250 = x93 & n4267;
  assign n11251 = x95 & n4270;
  assign n11252 = ~n11250 & ~n11251;
  assign n11253 = x94 & n4044;
  assign n11254 = n11252 & ~n11253;
  assign n11255 = ~n11249 & n11254;
  assign n11256 = n11255 ^ x38;
  assign n11371 = n11370 ^ n11256;
  assign n11246 = n11092 ^ n10990;
  assign n11247 = n11093 & n11246;
  assign n11248 = n11247 ^ n10990;
  assign n11372 = n11371 ^ n11248;
  assign n11238 = n3522 & n3763;
  assign n11239 = x96 & n3699;
  assign n11240 = x97 & n3526;
  assign n11241 = ~n11239 & ~n11240;
  assign n11242 = x98 & n3701;
  assign n11243 = n11241 & ~n11242;
  assign n11244 = ~n11238 & n11243;
  assign n11245 = n11244 ^ x35;
  assign n11373 = n11372 ^ n11245;
  assign n11235 = n11094 ^ n10979;
  assign n11236 = ~n11095 & ~n11235;
  assign n11237 = n11236 ^ n10979;
  assign n11374 = n11373 ^ n11237;
  assign n11227 = n3009 & n4323;
  assign n11228 = x100 & n3013;
  assign n11229 = x99 & n3181;
  assign n11230 = ~n11228 & ~n11229;
  assign n11231 = x101 & n3183;
  assign n11232 = n11230 & ~n11231;
  assign n11233 = ~n11227 & n11232;
  assign n11234 = n11233 ^ x32;
  assign n11375 = n11374 ^ n11234;
  assign n11224 = n11096 ^ n10968;
  assign n11225 = n11097 & n11224;
  assign n11226 = n11225 ^ n10968;
  assign n11376 = n11375 ^ n11226;
  assign n11216 = n2527 & n4912;
  assign n11217 = x103 & n2530;
  assign n11218 = x102 & n2690;
  assign n11219 = ~n11217 & ~n11218;
  assign n11220 = x104 & n2693;
  assign n11221 = n11219 & ~n11220;
  assign n11222 = ~n11216 & n11221;
  assign n11223 = n11222 ^ x29;
  assign n11377 = n11376 ^ n11223;
  assign n11213 = n11098 ^ n10957;
  assign n11214 = ~n11099 & ~n11213;
  assign n11215 = n11214 ^ n10957;
  assign n11378 = n11377 ^ n11215;
  assign n11205 = n2102 & n5578;
  assign n11206 = x105 & n2112;
  assign n11207 = x106 & n2105;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = x107 & n2381;
  assign n11210 = n11208 & ~n11209;
  assign n11211 = ~n11205 & n11210;
  assign n11212 = n11211 ^ x26;
  assign n11379 = n11378 ^ n11212;
  assign n11202 = n11100 ^ n10946;
  assign n11203 = n11101 & n11202;
  assign n11204 = n11203 ^ n10946;
  assign n11380 = n11379 ^ n11204;
  assign n11194 = n1746 & n6250;
  assign n11195 = x108 & n1871;
  assign n11196 = x109 & n1750;
  assign n11197 = ~n11195 & ~n11196;
  assign n11198 = x110 & n1873;
  assign n11199 = n11197 & ~n11198;
  assign n11200 = ~n11194 & n11199;
  assign n11201 = n11200 ^ x23;
  assign n11381 = n11380 ^ n11201;
  assign n11191 = n11102 ^ n10935;
  assign n11192 = ~n11103 & ~n11191;
  assign n11193 = n11192 ^ n10935;
  assign n11382 = n11381 ^ n11193;
  assign n11183 = n1404 & n6975;
  assign n11184 = x112 & n1408;
  assign n11185 = x111 & n1514;
  assign n11186 = ~n11184 & ~n11185;
  assign n11187 = x113 & n1517;
  assign n11188 = n11186 & ~n11187;
  assign n11189 = ~n11183 & n11188;
  assign n11190 = n11189 ^ x20;
  assign n11383 = n11382 ^ n11190;
  assign n11180 = n11104 ^ n10924;
  assign n11181 = n11105 & n11180;
  assign n11182 = n11181 ^ n10924;
  assign n11384 = n11383 ^ n11182;
  assign n11172 = n1098 & n7730;
  assign n11173 = x114 & n1198;
  assign n11174 = x115 & n1102;
  assign n11175 = ~n11173 & ~n11174;
  assign n11176 = x116 & n1201;
  assign n11177 = n11175 & ~n11176;
  assign n11178 = ~n11172 & n11177;
  assign n11179 = n11178 ^ x17;
  assign n11385 = n11384 ^ n11179;
  assign n11169 = n11106 ^ n10913;
  assign n11170 = ~n11107 & ~n11169;
  assign n11171 = n11170 ^ n10913;
  assign n11386 = n11385 ^ n11171;
  assign n11161 = n821 & n8542;
  assign n11162 = x117 & n898;
  assign n11163 = x119 & n901;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = x118 & n824;
  assign n11166 = n11164 & ~n11165;
  assign n11167 = ~n11161 & n11166;
  assign n11168 = n11167 ^ x14;
  assign n11387 = n11386 ^ n11168;
  assign n11158 = n11108 ^ n10902;
  assign n11159 = n11109 & n11158;
  assign n11160 = n11159 ^ n10902;
  assign n11388 = n11387 ^ n11160;
  assign n11150 = n596 & n9387;
  assign n11151 = x120 & n673;
  assign n11152 = x121 & n601;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = x122 & n676;
  assign n11155 = n11153 & ~n11154;
  assign n11156 = ~n11150 & n11155;
  assign n11157 = n11156 ^ x11;
  assign n11389 = n11388 ^ n11157;
  assign n11147 = n11110 ^ n10891;
  assign n11148 = ~n11111 & ~n11147;
  assign n11149 = n11148 ^ n10891;
  assign n11390 = n11389 ^ n11149;
  assign n11139 = n399 & n10303;
  assign n11140 = x123 & n478;
  assign n11141 = x124 & n402;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = x125 & n470;
  assign n11144 = n11142 & ~n11143;
  assign n11145 = ~n11139 & n11144;
  assign n11146 = n11145 ^ x8;
  assign n11391 = n11390 ^ n11146;
  assign n11136 = n11112 ^ n10880;
  assign n11137 = n11113 & n11136;
  assign n11138 = n11137 ^ n10880;
  assign n11392 = n11391 ^ n11138;
  assign n11130 = n239 & ~n10281;
  assign n11131 = x127 & n242;
  assign n11132 = x126 & n249;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~n11130 & n11133;
  assign n11135 = n11134 ^ x5;
  assign n11393 = n11392 ^ n11135;
  assign n11127 = n11114 ^ n10874;
  assign n11128 = n11115 & ~n11127;
  assign n11129 = n11128 ^ n10877;
  assign n11394 = n11393 ^ n11129;
  assign n11124 = n11116 ^ n10863;
  assign n11125 = ~n11117 & ~n11124;
  assign n11126 = n11125 ^ n10866;
  assign n11395 = n11394 ^ n11126;
  assign n11121 = n11118 ^ n10851;
  assign n11122 = ~n11119 & ~n11121;
  assign n11123 = n11122 ^ n10851;
  assign n11396 = n11395 ^ n11123;
  assign n11640 = n1667 & n6626;
  assign n11641 = x82 & n6884;
  assign n11642 = x83 & n6630;
  assign n11643 = ~n11641 & ~n11642;
  assign n11644 = x84 & n6888;
  assign n11645 = n11643 & ~n11644;
  assign n11646 = ~n11640 & n11645;
  assign n11647 = n11646 ^ x50;
  assign n11630 = n1340 & n7395;
  assign n11631 = x80 & n7400;
  assign n11632 = x79 & n7650;
  assign n11633 = ~n11631 & ~n11632;
  assign n11634 = x81 & n7652;
  assign n11635 = n11633 & ~n11634;
  assign n11636 = ~n11630 & n11635;
  assign n11637 = n11636 ^ x53;
  assign n11620 = n1041 & n8171;
  assign n11621 = x76 & n8181;
  assign n11622 = x78 & n8732;
  assign n11623 = ~n11621 & ~n11622;
  assign n11624 = x77 & n8174;
  assign n11625 = n11623 & ~n11624;
  assign n11626 = ~n11620 & n11625;
  assign n11627 = n11626 ^ x56;
  assign n11617 = n11329 ^ n11303;
  assign n11618 = n11330 & n11617;
  assign n11619 = n11618 ^ n11313;
  assign n11628 = n11627 ^ n11619;
  assign n11607 = n789 & n9002;
  assign n11608 = x73 & n9012;
  assign n11609 = x74 & n9005;
  assign n11610 = ~n11608 & ~n11609;
  assign n11611 = x75 & n9557;
  assign n11612 = n11610 & ~n11611;
  assign n11613 = ~n11607 & n11612;
  assign n11614 = n11613 ^ x59;
  assign n11597 = n11328 ^ x2;
  assign n11601 = n11316 ^ x2;
  assign n11602 = n11597 & n11601;
  assign n11603 = n11602 ^ x2;
  assign n11598 = n11317 ^ x2;
  assign n11599 = ~n11597 & n11598;
  assign n11600 = n11599 ^ x2;
  assign n11604 = n11603 ^ n11600;
  assign n11605 = ~x62 & n11604;
  assign n11606 = n11605 ^ n11603;
  assign n11615 = n11614 ^ n11606;
  assign n11589 = n575 & n9878;
  assign n11590 = x70 & n9888;
  assign n11591 = x72 & n10501;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = x71 & n9881;
  assign n11594 = n11592 & ~n11593;
  assign n11595 = ~n11589 & n11594;
  assign n11584 = x63 & x69;
  assign n11581 = x69 ^ x68;
  assign n11582 = ~x63 & n11581;
  assign n11583 = n11582 ^ x68;
  assign n11585 = n11584 ^ n11583;
  assign n11586 = ~x62 & ~n11585;
  assign n11587 = n11586 ^ n11583;
  assign n11588 = n11587 ^ x2;
  assign n11596 = n11595 ^ n11588;
  assign n11616 = n11615 ^ n11596;
  assign n11629 = n11628 ^ n11616;
  assign n11638 = n11637 ^ n11629;
  assign n11578 = n11331 ^ n11295;
  assign n11579 = n11340 & ~n11578;
  assign n11580 = n11579 ^ n11339;
  assign n11639 = n11638 ^ n11580;
  assign n11648 = n11647 ^ n11639;
  assign n11575 = n11349 ^ n11292;
  assign n11576 = ~n11350 & n11575;
  assign n11577 = n11576 ^ n11292;
  assign n11649 = n11648 ^ n11577;
  assign n11572 = n11362 ^ n11351;
  assign n11573 = ~n11363 & ~n11572;
  assign n11574 = n11573 ^ n11354;
  assign n11650 = n11649 ^ n11574;
  assign n11564 = n2039 & n5942;
  assign n11565 = x85 & n6186;
  assign n11566 = x87 & n6406;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = x86 & n5947;
  assign n11569 = n11567 & ~n11568;
  assign n11570 = ~n11564 & n11569;
  assign n11571 = n11570 ^ x47;
  assign n11651 = n11650 ^ n11571;
  assign n11556 = n2448 & n5262;
  assign n11557 = x88 & n5488;
  assign n11558 = x89 & n5266;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = x90 & n5491;
  assign n11561 = n11559 & ~n11560;
  assign n11562 = ~n11556 & n11561;
  assign n11563 = n11562 ^ x44;
  assign n11652 = n11651 ^ n11563;
  assign n11553 = n11364 ^ n11281;
  assign n11554 = n11365 & n11553;
  assign n11555 = n11554 ^ n11281;
  assign n11653 = n11652 ^ n11555;
  assign n11545 = n2901 & n4643;
  assign n11546 = x91 & n4653;
  assign n11547 = x93 & n5046;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = x92 & n4646;
  assign n11550 = n11548 & ~n11549;
  assign n11551 = ~n11545 & n11550;
  assign n11552 = n11551 ^ x41;
  assign n11654 = n11653 ^ n11552;
  assign n11542 = n11366 ^ n11270;
  assign n11543 = ~n11367 & ~n11542;
  assign n11544 = n11543 ^ n11270;
  assign n11655 = n11654 ^ n11544;
  assign n11534 = n3403 & n4040;
  assign n11535 = x94 & n4267;
  assign n11536 = x95 & n4044;
  assign n11537 = ~n11535 & ~n11536;
  assign n11538 = x96 & n4270;
  assign n11539 = n11537 & ~n11538;
  assign n11540 = ~n11534 & n11539;
  assign n11541 = n11540 ^ x38;
  assign n11656 = n11655 ^ n11541;
  assign n11531 = n11368 ^ n11259;
  assign n11532 = n11369 & n11531;
  assign n11533 = n11532 ^ n11259;
  assign n11657 = n11656 ^ n11533;
  assign n11523 = n3522 & n3943;
  assign n11524 = x97 & n3699;
  assign n11525 = x98 & n3526;
  assign n11526 = ~n11524 & ~n11525;
  assign n11527 = x99 & n3701;
  assign n11528 = n11526 & ~n11527;
  assign n11529 = ~n11523 & n11528;
  assign n11530 = n11529 ^ x35;
  assign n11658 = n11657 ^ n11530;
  assign n11520 = n11370 ^ n11248;
  assign n11521 = ~n11371 & ~n11520;
  assign n11522 = n11521 ^ n11248;
  assign n11659 = n11658 ^ n11522;
  assign n11512 = n3009 & n4509;
  assign n11513 = x100 & n3181;
  assign n11514 = x102 & n3183;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = x101 & n3013;
  assign n11517 = n11515 & ~n11516;
  assign n11518 = ~n11512 & n11517;
  assign n11519 = n11518 ^ x32;
  assign n11660 = n11659 ^ n11519;
  assign n11509 = n11372 ^ n11237;
  assign n11510 = n11373 & n11509;
  assign n11511 = n11510 ^ n11237;
  assign n11661 = n11660 ^ n11511;
  assign n11501 = n2527 & n5117;
  assign n11502 = x103 & n2690;
  assign n11503 = x104 & n2530;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = x105 & n2693;
  assign n11506 = n11504 & ~n11505;
  assign n11507 = ~n11501 & n11506;
  assign n11508 = n11507 ^ x29;
  assign n11662 = n11661 ^ n11508;
  assign n11498 = n11374 ^ n11226;
  assign n11499 = ~n11375 & ~n11498;
  assign n11500 = n11499 ^ n11226;
  assign n11663 = n11662 ^ n11500;
  assign n11490 = n2102 & n5792;
  assign n11491 = x106 & n2112;
  assign n11492 = x107 & n2105;
  assign n11493 = ~n11491 & ~n11492;
  assign n11494 = x108 & n2381;
  assign n11495 = n11493 & ~n11494;
  assign n11496 = ~n11490 & n11495;
  assign n11497 = n11496 ^ x26;
  assign n11664 = n11663 ^ n11497;
  assign n11487 = n11376 ^ n11215;
  assign n11488 = n11377 & n11487;
  assign n11489 = n11488 ^ n11215;
  assign n11665 = n11664 ^ n11489;
  assign n11479 = n1746 & n6478;
  assign n11480 = x109 & n1871;
  assign n11481 = x110 & n1750;
  assign n11482 = ~n11480 & ~n11481;
  assign n11483 = x111 & n1873;
  assign n11484 = n11482 & ~n11483;
  assign n11485 = ~n11479 & n11484;
  assign n11486 = n11485 ^ x23;
  assign n11666 = n11665 ^ n11486;
  assign n11476 = n11378 ^ n11204;
  assign n11477 = ~n11379 & ~n11476;
  assign n11478 = n11477 ^ n11204;
  assign n11667 = n11666 ^ n11478;
  assign n11468 = n1404 & n7220;
  assign n11469 = x112 & n1514;
  assign n11470 = x113 & n1408;
  assign n11471 = ~n11469 & ~n11470;
  assign n11472 = x114 & n1517;
  assign n11473 = n11471 & ~n11472;
  assign n11474 = ~n11468 & n11473;
  assign n11475 = n11474 ^ x20;
  assign n11668 = n11667 ^ n11475;
  assign n11465 = n11380 ^ n11193;
  assign n11466 = n11381 & n11465;
  assign n11467 = n11466 ^ n11193;
  assign n11669 = n11668 ^ n11467;
  assign n11457 = n1098 & n7987;
  assign n11458 = x115 & n1198;
  assign n11459 = x116 & n1102;
  assign n11460 = ~n11458 & ~n11459;
  assign n11461 = x117 & n1201;
  assign n11462 = n11460 & ~n11461;
  assign n11463 = ~n11457 & n11462;
  assign n11464 = n11463 ^ x17;
  assign n11670 = n11669 ^ n11464;
  assign n11454 = n11382 ^ n11182;
  assign n11455 = ~n11383 & ~n11454;
  assign n11456 = n11455 ^ n11182;
  assign n11671 = n11670 ^ n11456;
  assign n11446 = n821 & n8820;
  assign n11447 = x118 & n898;
  assign n11448 = x120 & n901;
  assign n11449 = ~n11447 & ~n11448;
  assign n11450 = x119 & n824;
  assign n11451 = n11449 & ~n11450;
  assign n11452 = ~n11446 & n11451;
  assign n11453 = n11452 ^ x14;
  assign n11672 = n11671 ^ n11453;
  assign n11443 = n11384 ^ n11171;
  assign n11444 = n11385 & n11443;
  assign n11445 = n11444 ^ n11171;
  assign n11673 = n11672 ^ n11445;
  assign n11435 = n596 & n9691;
  assign n11436 = x121 & n673;
  assign n11437 = x122 & n601;
  assign n11438 = ~n11436 & ~n11437;
  assign n11439 = x123 & n676;
  assign n11440 = n11438 & ~n11439;
  assign n11441 = ~n11435 & n11440;
  assign n11442 = n11441 ^ x11;
  assign n11674 = n11673 ^ n11442;
  assign n11432 = n11386 ^ n11160;
  assign n11433 = ~n11387 & ~n11432;
  assign n11434 = n11433 ^ n11160;
  assign n11675 = n11674 ^ n11434;
  assign n11424 = n399 & ~n10570;
  assign n11425 = x124 & n478;
  assign n11426 = x125 & n402;
  assign n11427 = ~n11425 & ~n11426;
  assign n11428 = x126 & n470;
  assign n11429 = n11427 & ~n11428;
  assign n11430 = ~n11424 & n11429;
  assign n11431 = n11430 ^ x8;
  assign n11676 = n11675 ^ n11431;
  assign n11421 = n11388 ^ n11149;
  assign n11422 = n11389 & n11421;
  assign n11423 = n11422 ^ n11149;
  assign n11677 = n11676 ^ n11423;
  assign n11406 = x127 & n183;
  assign n11407 = ~x5 & ~n11406;
  assign n11408 = n11407 ^ x4;
  assign n11409 = x127 & ~n10278;
  assign n11410 = n178 & n11409;
  assign n11411 = n11410 ^ n11407;
  assign n11412 = ~n11407 & n11411;
  assign n11413 = n11412 ^ n11407;
  assign n11414 = x127 & n248;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = n11415 ^ n11412;
  assign n11417 = n11416 ^ n11407;
  assign n11418 = n11417 ^ n11410;
  assign n11419 = ~n11408 & n11418;
  assign n11420 = n11419 ^ x4;
  assign n11678 = n11677 ^ n11420;
  assign n11403 = n11390 ^ n11138;
  assign n11404 = ~n11391 & ~n11403;
  assign n11405 = n11404 ^ n11138;
  assign n11679 = n11678 ^ n11405;
  assign n11400 = n11392 ^ n11129;
  assign n11401 = n11393 & ~n11400;
  assign n11402 = n11401 ^ n11129;
  assign n11680 = n11679 ^ n11402;
  assign n11397 = n11126 ^ n11123;
  assign n11398 = ~n11395 & ~n11397;
  assign n11399 = n11398 ^ n11123;
  assign n11681 = n11680 ^ n11399;
  assign n11941 = ~n11402 & n11677;
  assign n11942 = ~n11405 & ~n11420;
  assign n11948 = ~n11941 & n11942;
  assign n11944 = n11402 & ~n11677;
  assign n11945 = n11405 & n11420;
  assign n11949 = n11944 & ~n11945;
  assign n11950 = ~n11948 & ~n11949;
  assign n11943 = n11941 & ~n11942;
  assign n11946 = ~n11944 & n11945;
  assign n11947 = ~n11943 & ~n11946;
  assign n11951 = n11950 ^ n11947;
  assign n11952 = ~n11399 & n11951;
  assign n11953 = n11952 ^ n11950;
  assign n11954 = n11405 ^ n11402;
  assign n11955 = n11677 ^ n11405;
  assign n11956 = ~n11678 & ~n11955;
  assign n11957 = n11954 & n11956;
  assign n11958 = n11953 & ~n11957;
  assign n11899 = n1149 & n8171;
  assign n11900 = x77 & n8181;
  assign n11901 = x78 & n8174;
  assign n11902 = ~n11900 & ~n11901;
  assign n11903 = x79 & n8732;
  assign n11904 = n11902 & ~n11903;
  assign n11905 = ~n11899 & n11904;
  assign n11906 = n11905 ^ x56;
  assign n11896 = n11619 ^ n11616;
  assign n11897 = ~n11628 & n11896;
  assign n11898 = n11897 ^ n11627;
  assign n11907 = n11906 ^ n11898;
  assign n11890 = x5 ^ x2;
  assign n11887 = n11584 ^ x70;
  assign n11888 = ~n10177 & n11887;
  assign n11889 = n11888 ^ x70;
  assign n11891 = n11890 ^ n11889;
  assign n11877 = n11595 ^ x2;
  assign n11881 = n11583 ^ x2;
  assign n11882 = n11877 & n11881;
  assign n11883 = n11882 ^ x2;
  assign n11878 = n11584 ^ x2;
  assign n11879 = ~n11877 & n11878;
  assign n11880 = n11879 ^ x2;
  assign n11884 = n11883 ^ n11880;
  assign n11885 = ~x62 & n11884;
  assign n11886 = n11885 ^ n11883;
  assign n11892 = n11891 ^ n11886;
  assign n11869 = ~n653 & n9878;
  assign n11870 = x71 & n9888;
  assign n11871 = x73 & n10501;
  assign n11872 = ~n11870 & ~n11871;
  assign n11873 = x72 & n9881;
  assign n11874 = n11872 & ~n11873;
  assign n11875 = ~n11869 & n11874;
  assign n11876 = n11875 ^ x62;
  assign n11893 = n11892 ^ n11876;
  assign n11861 = n870 & n9002;
  assign n11862 = x74 & n9012;
  assign n11863 = x75 & n9005;
  assign n11864 = ~n11862 & ~n11863;
  assign n11865 = x76 & n9557;
  assign n11866 = n11864 & ~n11865;
  assign n11867 = ~n11861 & n11866;
  assign n11868 = n11867 ^ x59;
  assign n11894 = n11893 ^ n11868;
  assign n11858 = n11606 ^ n11596;
  assign n11859 = ~n11615 & ~n11858;
  assign n11860 = n11859 ^ n11614;
  assign n11895 = n11894 ^ n11860;
  assign n11908 = n11907 ^ n11895;
  assign n11850 = n1454 & n7395;
  assign n11851 = x80 & n7650;
  assign n11852 = x81 & n7400;
  assign n11853 = ~n11851 & ~n11852;
  assign n11854 = x82 & n7652;
  assign n11855 = n11853 & ~n11854;
  assign n11856 = ~n11850 & n11855;
  assign n11857 = n11856 ^ x53;
  assign n11909 = n11908 ^ n11857;
  assign n11847 = n11629 ^ n11580;
  assign n11848 = ~n11638 & n11847;
  assign n11849 = n11848 ^ n11637;
  assign n11910 = n11909 ^ n11849;
  assign n11839 = n1801 & n6626;
  assign n11840 = x83 & n6884;
  assign n11841 = x85 & n6888;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = x84 & n6630;
  assign n11844 = n11842 & ~n11843;
  assign n11845 = ~n11839 & n11844;
  assign n11846 = n11845 ^ x50;
  assign n11911 = n11910 ^ n11846;
  assign n11836 = n11647 ^ n11577;
  assign n11837 = n11648 & n11836;
  assign n11838 = n11837 ^ n11577;
  assign n11912 = n11911 ^ n11838;
  assign n11833 = n11649 ^ n11571;
  assign n11834 = n11650 & n11833;
  assign n11835 = n11834 ^ n11574;
  assign n11913 = n11912 ^ n11835;
  assign n11825 = n2176 & n5942;
  assign n11826 = x86 & n6186;
  assign n11827 = x88 & n6406;
  assign n11828 = ~n11826 & ~n11827;
  assign n11829 = x87 & n5947;
  assign n11830 = n11828 & ~n11829;
  assign n11831 = ~n11825 & n11830;
  assign n11832 = n11831 ^ x47;
  assign n11914 = n11913 ^ n11832;
  assign n11817 = n2607 & n5262;
  assign n11818 = x89 & n5488;
  assign n11819 = x91 & n5491;
  assign n11820 = ~n11818 & ~n11819;
  assign n11821 = x90 & n5266;
  assign n11822 = n11820 & ~n11821;
  assign n11823 = ~n11817 & n11822;
  assign n11824 = n11823 ^ x44;
  assign n11915 = n11914 ^ n11824;
  assign n11814 = n11651 ^ n11555;
  assign n11815 = ~n11652 & ~n11814;
  assign n11816 = n11815 ^ n11555;
  assign n11916 = n11915 ^ n11816;
  assign n11806 = n3078 & n4643;
  assign n11807 = x92 & n4653;
  assign n11808 = x93 & n4646;
  assign n11809 = ~n11807 & ~n11808;
  assign n11810 = x94 & n5046;
  assign n11811 = n11809 & ~n11810;
  assign n11812 = ~n11806 & n11811;
  assign n11813 = n11812 ^ x41;
  assign n11917 = n11916 ^ n11813;
  assign n11803 = n11653 ^ n11544;
  assign n11804 = n11654 & n11803;
  assign n11805 = n11804 ^ n11544;
  assign n11918 = n11917 ^ n11805;
  assign n11795 = n3585 & n4040;
  assign n11796 = x95 & n4267;
  assign n11797 = x97 & n4270;
  assign n11798 = ~n11796 & ~n11797;
  assign n11799 = x96 & n4044;
  assign n11800 = n11798 & ~n11799;
  assign n11801 = ~n11795 & n11800;
  assign n11802 = n11801 ^ x38;
  assign n11919 = n11918 ^ n11802;
  assign n11792 = n11655 ^ n11533;
  assign n11793 = ~n11656 & ~n11792;
  assign n11794 = n11793 ^ n11533;
  assign n11920 = n11919 ^ n11794;
  assign n11784 = n3522 & n4141;
  assign n11785 = x98 & n3699;
  assign n11786 = x99 & n3526;
  assign n11787 = ~n11785 & ~n11786;
  assign n11788 = x100 & n3701;
  assign n11789 = n11787 & ~n11788;
  assign n11790 = ~n11784 & n11789;
  assign n11791 = n11790 ^ x35;
  assign n11921 = n11920 ^ n11791;
  assign n11781 = n11657 ^ n11522;
  assign n11782 = n11658 & n11781;
  assign n11783 = n11782 ^ n11522;
  assign n11922 = n11921 ^ n11783;
  assign n11773 = n3009 & n4718;
  assign n11774 = x101 & n3181;
  assign n11775 = x102 & n3013;
  assign n11776 = ~n11774 & ~n11775;
  assign n11777 = x103 & n3183;
  assign n11778 = n11776 & ~n11777;
  assign n11779 = ~n11773 & n11778;
  assign n11780 = n11779 ^ x32;
  assign n11923 = n11922 ^ n11780;
  assign n11770 = n11659 ^ n11511;
  assign n11771 = ~n11660 & ~n11770;
  assign n11772 = n11771 ^ n11511;
  assign n11924 = n11923 ^ n11772;
  assign n11762 = n2527 & n5351;
  assign n11763 = x104 & n2690;
  assign n11764 = x105 & n2530;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = x106 & n2693;
  assign n11767 = n11765 & ~n11766;
  assign n11768 = ~n11762 & n11767;
  assign n11769 = n11768 ^ x29;
  assign n11925 = n11924 ^ n11769;
  assign n11759 = n11661 ^ n11500;
  assign n11760 = n11662 & n11759;
  assign n11761 = n11760 ^ n11500;
  assign n11926 = n11925 ^ n11761;
  assign n11751 = n2102 & n6026;
  assign n11752 = x107 & n2112;
  assign n11753 = x108 & n2105;
  assign n11754 = ~n11752 & ~n11753;
  assign n11755 = x109 & n2381;
  assign n11756 = n11754 & ~n11755;
  assign n11757 = ~n11751 & n11756;
  assign n11758 = n11757 ^ x26;
  assign n11927 = n11926 ^ n11758;
  assign n11748 = n11663 ^ n11489;
  assign n11749 = ~n11664 & ~n11748;
  assign n11750 = n11749 ^ n11489;
  assign n11928 = n11927 ^ n11750;
  assign n11740 = n1746 & n6728;
  assign n11741 = x111 & n1750;
  assign n11742 = x110 & n1871;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = x112 & n1873;
  assign n11745 = n11743 & ~n11744;
  assign n11746 = ~n11740 & n11745;
  assign n11747 = n11746 ^ x23;
  assign n11929 = n11928 ^ n11747;
  assign n11737 = n11665 ^ n11478;
  assign n11738 = n11666 & n11737;
  assign n11739 = n11738 ^ n11478;
  assign n11930 = n11929 ^ n11739;
  assign n11729 = n1404 & n7481;
  assign n11730 = x113 & n1514;
  assign n11731 = x114 & n1408;
  assign n11732 = ~n11730 & ~n11731;
  assign n11733 = x115 & n1517;
  assign n11734 = n11732 & ~n11733;
  assign n11735 = ~n11729 & n11734;
  assign n11736 = n11735 ^ x20;
  assign n11931 = n11930 ^ n11736;
  assign n11726 = n11667 ^ n11467;
  assign n11727 = ~n11668 & ~n11726;
  assign n11728 = n11727 ^ n11467;
  assign n11932 = n11931 ^ n11728;
  assign n11718 = n1098 & n8265;
  assign n11719 = x116 & n1198;
  assign n11720 = x117 & n1102;
  assign n11721 = ~n11719 & ~n11720;
  assign n11722 = x118 & n1201;
  assign n11723 = n11721 & ~n11722;
  assign n11724 = ~n11718 & n11723;
  assign n11725 = n11724 ^ x17;
  assign n11933 = n11932 ^ n11725;
  assign n11715 = n11669 ^ n11456;
  assign n11716 = n11670 & n11715;
  assign n11717 = n11716 ^ n11456;
  assign n11934 = n11933 ^ n11717;
  assign n11707 = n821 & n9094;
  assign n11708 = x120 & n824;
  assign n11709 = x119 & n898;
  assign n11710 = ~n11708 & ~n11709;
  assign n11711 = x121 & n901;
  assign n11712 = n11710 & ~n11711;
  assign n11713 = ~n11707 & n11712;
  assign n11714 = n11713 ^ x14;
  assign n11935 = n11934 ^ n11714;
  assign n11704 = n11671 ^ n11445;
  assign n11705 = ~n11672 & ~n11704;
  assign n11706 = n11705 ^ n11445;
  assign n11936 = n11935 ^ n11706;
  assign n11696 = n596 & n9999;
  assign n11697 = x122 & n673;
  assign n11698 = x123 & n601;
  assign n11699 = ~n11697 & ~n11698;
  assign n11700 = x124 & n676;
  assign n11701 = n11699 & ~n11700;
  assign n11702 = ~n11696 & n11701;
  assign n11703 = n11702 ^ x11;
  assign n11937 = n11936 ^ n11703;
  assign n11693 = n11673 ^ n11434;
  assign n11694 = n11674 & n11693;
  assign n11695 = n11694 ^ n11434;
  assign n11938 = n11937 ^ n11695;
  assign n11685 = n399 & ~n10855;
  assign n11686 = x125 & n478;
  assign n11687 = x126 & n402;
  assign n11688 = ~n11686 & ~n11687;
  assign n11689 = x127 & n470;
  assign n11690 = n11688 & ~n11689;
  assign n11691 = ~n11685 & n11690;
  assign n11692 = n11691 ^ x8;
  assign n11939 = n11938 ^ n11692;
  assign n11682 = n11675 ^ n11423;
  assign n11683 = ~n11676 & ~n11682;
  assign n11684 = n11683 ^ n11423;
  assign n11940 = n11939 ^ n11684;
  assign n11959 = n11958 ^ n11940;
  assign n12213 = ~n11940 & ~n11944;
  assign n12214 = n11399 & ~n12213;
  assign n12215 = n11940 & ~n11941;
  assign n12216 = ~n11942 & ~n12215;
  assign n12217 = ~n12214 & n12216;
  assign n12218 = ~n11940 & n11945;
  assign n12219 = ~n12217 & ~n12218;
  assign n12220 = n11399 & ~n11941;
  assign n12221 = ~n11946 & ~n12213;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = n12219 & ~n12222;
  assign n12178 = n2755 & n5262;
  assign n12179 = x90 & n5488;
  assign n12180 = x92 & n5491;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = x91 & n5266;
  assign n12183 = n12181 & ~n12182;
  assign n12184 = ~n12178 & n12183;
  assign n12185 = n12184 ^ x44;
  assign n12168 = n2310 & n5942;
  assign n12169 = x87 & n6186;
  assign n12170 = x88 & n5947;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = x89 & n6406;
  assign n12173 = n12171 & ~n12172;
  assign n12174 = ~n12168 & n12173;
  assign n12175 = n12174 ^ x47;
  assign n12158 = n1920 & n6626;
  assign n12159 = x84 & n6884;
  assign n12160 = x86 & n6888;
  assign n12161 = ~n12159 & ~n12160;
  assign n12162 = x85 & n6630;
  assign n12163 = n12161 & ~n12162;
  assign n12164 = ~n12158 & n12163;
  assign n12165 = n12164 ^ x50;
  assign n12148 = n1560 & n7395;
  assign n12149 = x81 & n7650;
  assign n12150 = x82 & n7400;
  assign n12151 = ~n12149 & ~n12150;
  assign n12152 = x83 & n7652;
  assign n12153 = n12151 & ~n12152;
  assign n12154 = ~n12148 & n12153;
  assign n12155 = n12154 ^ x53;
  assign n12136 = n956 & n9002;
  assign n12137 = x75 & n9012;
  assign n12138 = x77 & n9557;
  assign n12139 = ~n12137 & ~n12138;
  assign n12140 = x76 & n9005;
  assign n12141 = n12139 & ~n12140;
  assign n12142 = ~n12136 & n12141;
  assign n12143 = n12142 ^ x59;
  assign n12127 = ~n721 & n9878;
  assign n12128 = x73 & n9881;
  assign n12129 = x72 & n9888;
  assign n12130 = ~n12128 & ~n12129;
  assign n12131 = x74 & n10501;
  assign n12132 = n12130 & ~n12131;
  assign n12133 = ~n12127 & n12132;
  assign n12134 = n12133 ^ x62;
  assign n12122 = x71 & n10177;
  assign n12123 = x62 & x63;
  assign n12124 = x70 & n12123;
  assign n12125 = ~n12122 & ~n12124;
  assign n12119 = n11889 ^ x5;
  assign n12120 = n11890 & n12119;
  assign n12121 = n12120 ^ x2;
  assign n12126 = n12125 ^ n12121;
  assign n12135 = n12134 ^ n12126;
  assign n12144 = n12143 ^ n12135;
  assign n12116 = n11891 ^ n11876;
  assign n12117 = n11892 & n12116;
  assign n12118 = n12117 ^ n11886;
  assign n12145 = n12144 ^ n12118;
  assign n12108 = n1242 & n8171;
  assign n12109 = x78 & n8181;
  assign n12110 = x79 & n8174;
  assign n12111 = ~n12109 & ~n12110;
  assign n12112 = x80 & n8732;
  assign n12113 = n12111 & ~n12112;
  assign n12114 = ~n12108 & n12113;
  assign n12115 = n12114 ^ x56;
  assign n12146 = n12145 ^ n12115;
  assign n12105 = n11893 ^ n11860;
  assign n12106 = ~n11894 & n12105;
  assign n12107 = n12106 ^ n11860;
  assign n12147 = n12146 ^ n12107;
  assign n12156 = n12155 ^ n12147;
  assign n12102 = n11906 ^ n11895;
  assign n12103 = n11907 & ~n12102;
  assign n12104 = n12103 ^ n11898;
  assign n12157 = n12156 ^ n12104;
  assign n12166 = n12165 ^ n12157;
  assign n12099 = n11857 ^ n11849;
  assign n12100 = n11909 & ~n12099;
  assign n12101 = n12100 ^ n11908;
  assign n12167 = n12166 ^ n12101;
  assign n12176 = n12175 ^ n12167;
  assign n12096 = n11910 ^ n11838;
  assign n12097 = ~n11911 & n12096;
  assign n12098 = n12097 ^ n11838;
  assign n12177 = n12176 ^ n12098;
  assign n12186 = n12185 ^ n12177;
  assign n12093 = n11912 ^ n11832;
  assign n12094 = ~n11913 & ~n12093;
  assign n12095 = n12094 ^ n11835;
  assign n12187 = n12186 ^ n12095;
  assign n12085 = n3247 & n4643;
  assign n12086 = x93 & n4653;
  assign n12087 = x95 & n5046;
  assign n12088 = ~n12086 & ~n12087;
  assign n12089 = x94 & n4646;
  assign n12090 = n12088 & ~n12089;
  assign n12091 = ~n12085 & n12090;
  assign n12092 = n12091 ^ x41;
  assign n12188 = n12187 ^ n12092;
  assign n12082 = n11914 ^ n11816;
  assign n12083 = n11915 & n12082;
  assign n12084 = n12083 ^ n11816;
  assign n12189 = n12188 ^ n12084;
  assign n12074 = n3763 & n4040;
  assign n12075 = x96 & n4267;
  assign n12076 = x98 & n4270;
  assign n12077 = ~n12075 & ~n12076;
  assign n12078 = x97 & n4044;
  assign n12079 = n12077 & ~n12078;
  assign n12080 = ~n12074 & n12079;
  assign n12081 = n12080 ^ x38;
  assign n12190 = n12189 ^ n12081;
  assign n12071 = n11916 ^ n11805;
  assign n12072 = ~n11917 & ~n12071;
  assign n12073 = n12072 ^ n11805;
  assign n12191 = n12190 ^ n12073;
  assign n12063 = n3522 & n4323;
  assign n12064 = x99 & n3699;
  assign n12065 = x100 & n3526;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = x101 & n3701;
  assign n12068 = n12066 & ~n12067;
  assign n12069 = ~n12063 & n12068;
  assign n12070 = n12069 ^ x35;
  assign n12192 = n12191 ^ n12070;
  assign n12060 = n11918 ^ n11794;
  assign n12061 = n11919 & n12060;
  assign n12062 = n12061 ^ n11794;
  assign n12193 = n12192 ^ n12062;
  assign n12052 = n3009 & n4912;
  assign n12053 = x103 & n3013;
  assign n12054 = x102 & n3181;
  assign n12055 = ~n12053 & ~n12054;
  assign n12056 = x104 & n3183;
  assign n12057 = n12055 & ~n12056;
  assign n12058 = ~n12052 & n12057;
  assign n12059 = n12058 ^ x32;
  assign n12194 = n12193 ^ n12059;
  assign n12049 = n11920 ^ n11783;
  assign n12050 = ~n11921 & ~n12049;
  assign n12051 = n12050 ^ n11783;
  assign n12195 = n12194 ^ n12051;
  assign n12041 = n2527 & n5578;
  assign n12042 = x105 & n2690;
  assign n12043 = x106 & n2530;
  assign n12044 = ~n12042 & ~n12043;
  assign n12045 = x107 & n2693;
  assign n12046 = n12044 & ~n12045;
  assign n12047 = ~n12041 & n12046;
  assign n12048 = n12047 ^ x29;
  assign n12196 = n12195 ^ n12048;
  assign n12038 = n11922 ^ n11772;
  assign n12039 = n11923 & n12038;
  assign n12040 = n12039 ^ n11772;
  assign n12197 = n12196 ^ n12040;
  assign n12030 = n2102 & n6250;
  assign n12031 = x108 & n2112;
  assign n12032 = x109 & n2105;
  assign n12033 = ~n12031 & ~n12032;
  assign n12034 = x110 & n2381;
  assign n12035 = n12033 & ~n12034;
  assign n12036 = ~n12030 & n12035;
  assign n12037 = n12036 ^ x26;
  assign n12198 = n12197 ^ n12037;
  assign n12027 = n11924 ^ n11761;
  assign n12028 = ~n11925 & ~n12027;
  assign n12029 = n12028 ^ n11761;
  assign n12199 = n12198 ^ n12029;
  assign n12019 = n1746 & n6975;
  assign n12020 = x112 & n1750;
  assign n12021 = x111 & n1871;
  assign n12022 = ~n12020 & ~n12021;
  assign n12023 = x113 & n1873;
  assign n12024 = n12022 & ~n12023;
  assign n12025 = ~n12019 & n12024;
  assign n12026 = n12025 ^ x23;
  assign n12200 = n12199 ^ n12026;
  assign n12016 = n11926 ^ n11750;
  assign n12017 = n11927 & n12016;
  assign n12018 = n12017 ^ n11750;
  assign n12201 = n12200 ^ n12018;
  assign n12008 = n1404 & n7730;
  assign n12009 = x114 & n1514;
  assign n12010 = x115 & n1408;
  assign n12011 = ~n12009 & ~n12010;
  assign n12012 = x116 & n1517;
  assign n12013 = n12011 & ~n12012;
  assign n12014 = ~n12008 & n12013;
  assign n12015 = n12014 ^ x20;
  assign n12202 = n12201 ^ n12015;
  assign n12005 = n11928 ^ n11739;
  assign n12006 = ~n11929 & ~n12005;
  assign n12007 = n12006 ^ n11739;
  assign n12203 = n12202 ^ n12007;
  assign n11997 = n1098 & n8542;
  assign n11998 = x117 & n1198;
  assign n11999 = x118 & n1102;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = x119 & n1201;
  assign n12002 = n12000 & ~n12001;
  assign n12003 = ~n11997 & n12002;
  assign n12004 = n12003 ^ x17;
  assign n12204 = n12203 ^ n12004;
  assign n11994 = n11930 ^ n11728;
  assign n11995 = n11931 & n11994;
  assign n11996 = n11995 ^ n11728;
  assign n12205 = n12204 ^ n11996;
  assign n11986 = n821 & n9387;
  assign n11987 = x120 & n898;
  assign n11988 = x121 & n824;
  assign n11989 = ~n11987 & ~n11988;
  assign n11990 = x122 & n901;
  assign n11991 = n11989 & ~n11990;
  assign n11992 = ~n11986 & n11991;
  assign n11993 = n11992 ^ x14;
  assign n12206 = n12205 ^ n11993;
  assign n11983 = n11932 ^ n11717;
  assign n11984 = ~n11933 & ~n11983;
  assign n11985 = n11984 ^ n11717;
  assign n12207 = n12206 ^ n11985;
  assign n11975 = n596 & n10303;
  assign n11976 = x123 & n673;
  assign n11977 = x124 & n601;
  assign n11978 = ~n11976 & ~n11977;
  assign n11979 = x125 & n676;
  assign n11980 = n11978 & ~n11979;
  assign n11981 = ~n11975 & n11980;
  assign n11982 = n11981 ^ x11;
  assign n12208 = n12207 ^ n11982;
  assign n11972 = n11934 ^ n11706;
  assign n11973 = n11935 & n11972;
  assign n11974 = n11973 ^ n11706;
  assign n12209 = n12208 ^ n11974;
  assign n11966 = n399 & ~n10281;
  assign n11967 = x126 & n478;
  assign n11968 = x127 & n402;
  assign n11969 = ~n11967 & ~n11968;
  assign n11970 = ~n11966 & n11969;
  assign n11971 = n11970 ^ x8;
  assign n12210 = n12209 ^ n11971;
  assign n11963 = n11936 ^ n11695;
  assign n11964 = ~n11937 & ~n11963;
  assign n11965 = n11964 ^ n11695;
  assign n12211 = n12210 ^ n11965;
  assign n11960 = n11938 ^ n11684;
  assign n11961 = n11939 & n11960;
  assign n11962 = n11961 ^ n11684;
  assign n12212 = n12211 ^ n11962;
  assign n12224 = n12223 ^ n12212;
  assign n12455 = n3403 & n4643;
  assign n12456 = x94 & n4653;
  assign n12457 = x95 & n4646;
  assign n12458 = ~n12456 & ~n12457;
  assign n12459 = x96 & n5046;
  assign n12460 = n12458 & ~n12459;
  assign n12461 = ~n12455 & n12460;
  assign n12462 = n12461 ^ x41;
  assign n12445 = n2901 & n5262;
  assign n12446 = x91 & n5488;
  assign n12447 = x92 & n5266;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = x93 & n5491;
  assign n12450 = n12448 & ~n12449;
  assign n12451 = ~n12445 & n12450;
  assign n12452 = n12451 ^ x44;
  assign n12435 = n2448 & n5942;
  assign n12436 = x88 & n6186;
  assign n12437 = x90 & n6406;
  assign n12438 = ~n12436 & ~n12437;
  assign n12439 = x89 & n5947;
  assign n12440 = n12438 & ~n12439;
  assign n12441 = ~n12435 & n12440;
  assign n12442 = n12441 ^ x47;
  assign n12432 = n12165 ^ n12101;
  assign n12433 = ~n12166 & n12432;
  assign n12434 = n12433 ^ n12101;
  assign n12443 = n12442 ^ n12434;
  assign n12422 = n2039 & n6626;
  assign n12423 = x85 & n6884;
  assign n12424 = x87 & n6888;
  assign n12425 = ~n12423 & ~n12424;
  assign n12426 = x86 & n6630;
  assign n12427 = n12425 & ~n12426;
  assign n12428 = ~n12422 & n12427;
  assign n12429 = n12428 ^ x50;
  assign n12412 = n1667 & n7395;
  assign n12413 = x82 & n7650;
  assign n12414 = x83 & n7400;
  assign n12415 = ~n12413 & ~n12414;
  assign n12416 = x84 & n7652;
  assign n12417 = n12415 & ~n12416;
  assign n12418 = ~n12412 & n12417;
  assign n12419 = n12418 ^ x53;
  assign n12400 = n1041 & n9002;
  assign n12401 = x76 & n9012;
  assign n12402 = x77 & n9005;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = x78 & n9557;
  assign n12405 = n12403 & ~n12404;
  assign n12406 = ~n12400 & n12405;
  assign n12407 = n12406 ^ x59;
  assign n12392 = n789 & n9878;
  assign n12393 = x73 & n9888;
  assign n12394 = x74 & n9881;
  assign n12395 = ~n12393 & ~n12394;
  assign n12396 = x75 & n10501;
  assign n12397 = n12395 & ~n12396;
  assign n12398 = ~n12392 & n12397;
  assign n12399 = n12398 ^ x62;
  assign n12408 = n12407 ^ n12399;
  assign n12388 = n12134 ^ n12121;
  assign n12389 = n12126 & n12388;
  assign n12390 = n12389 ^ n12134;
  assign n12379 = x72 ^ x71;
  assign n12380 = n12379 ^ x63;
  assign n12381 = n12380 ^ n12379;
  assign n12382 = n12379 ^ n377;
  assign n12383 = n12382 ^ n12379;
  assign n12384 = n12381 & n12383;
  assign n12385 = n12384 ^ n12379;
  assign n12386 = ~n10177 & n12385;
  assign n12387 = n12386 ^ n12379;
  assign n12391 = n12390 ^ n12387;
  assign n12409 = n12408 ^ n12391;
  assign n12371 = n1340 & n8171;
  assign n12372 = x79 & n8181;
  assign n12373 = x81 & n8732;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = x80 & n8174;
  assign n12376 = n12374 & ~n12375;
  assign n12377 = ~n12371 & n12376;
  assign n12378 = n12377 ^ x56;
  assign n12410 = n12409 ^ n12378;
  assign n12368 = n12143 ^ n12118;
  assign n12369 = n12144 & ~n12368;
  assign n12370 = n12369 ^ n12118;
  assign n12411 = n12410 ^ n12370;
  assign n12420 = n12419 ^ n12411;
  assign n12365 = n12145 ^ n12107;
  assign n12366 = ~n12146 & n12365;
  assign n12367 = n12366 ^ n12107;
  assign n12421 = n12420 ^ n12367;
  assign n12430 = n12429 ^ n12421;
  assign n12362 = n12155 ^ n12104;
  assign n12363 = ~n12156 & n12362;
  assign n12364 = n12363 ^ n12104;
  assign n12431 = n12430 ^ n12364;
  assign n12444 = n12443 ^ n12431;
  assign n12453 = n12452 ^ n12444;
  assign n12359 = n12167 ^ n12098;
  assign n12360 = n12176 & ~n12359;
  assign n12361 = n12360 ^ n12175;
  assign n12454 = n12453 ^ n12361;
  assign n12463 = n12462 ^ n12454;
  assign n12356 = n12185 ^ n12095;
  assign n12357 = ~n12186 & ~n12356;
  assign n12358 = n12357 ^ n12095;
  assign n12464 = n12463 ^ n12358;
  assign n12348 = n3943 & n4040;
  assign n12349 = x97 & n4267;
  assign n12350 = x99 & n4270;
  assign n12351 = ~n12349 & ~n12350;
  assign n12352 = x98 & n4044;
  assign n12353 = n12351 & ~n12352;
  assign n12354 = ~n12348 & n12353;
  assign n12355 = n12354 ^ x38;
  assign n12465 = n12464 ^ n12355;
  assign n12345 = n12187 ^ n12084;
  assign n12346 = n12188 & n12345;
  assign n12347 = n12346 ^ n12084;
  assign n12466 = n12465 ^ n12347;
  assign n12337 = n3522 & n4509;
  assign n12338 = x100 & n3699;
  assign n12339 = x102 & n3701;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = x101 & n3526;
  assign n12342 = n12340 & ~n12341;
  assign n12343 = ~n12337 & n12342;
  assign n12344 = n12343 ^ x35;
  assign n12467 = n12466 ^ n12344;
  assign n12334 = n12189 ^ n12073;
  assign n12335 = ~n12190 & ~n12334;
  assign n12336 = n12335 ^ n12073;
  assign n12468 = n12467 ^ n12336;
  assign n12326 = n3009 & n5117;
  assign n12327 = x103 & n3181;
  assign n12328 = x104 & n3013;
  assign n12329 = ~n12327 & ~n12328;
  assign n12330 = x105 & n3183;
  assign n12331 = n12329 & ~n12330;
  assign n12332 = ~n12326 & n12331;
  assign n12333 = n12332 ^ x32;
  assign n12469 = n12468 ^ n12333;
  assign n12323 = n12191 ^ n12062;
  assign n12324 = n12192 & n12323;
  assign n12325 = n12324 ^ n12062;
  assign n12470 = n12469 ^ n12325;
  assign n12315 = n2527 & n5792;
  assign n12316 = x107 & n2530;
  assign n12317 = x106 & n2690;
  assign n12318 = ~n12316 & ~n12317;
  assign n12319 = x108 & n2693;
  assign n12320 = n12318 & ~n12319;
  assign n12321 = ~n12315 & n12320;
  assign n12322 = n12321 ^ x29;
  assign n12471 = n12470 ^ n12322;
  assign n12312 = n12193 ^ n12051;
  assign n12313 = ~n12194 & ~n12312;
  assign n12314 = n12313 ^ n12051;
  assign n12472 = n12471 ^ n12314;
  assign n12304 = n2102 & n6478;
  assign n12305 = x109 & n2112;
  assign n12306 = x111 & n2381;
  assign n12307 = ~n12305 & ~n12306;
  assign n12308 = x110 & n2105;
  assign n12309 = n12307 & ~n12308;
  assign n12310 = ~n12304 & n12309;
  assign n12311 = n12310 ^ x26;
  assign n12473 = n12472 ^ n12311;
  assign n12301 = n12195 ^ n12040;
  assign n12302 = n12196 & n12301;
  assign n12303 = n12302 ^ n12040;
  assign n12474 = n12473 ^ n12303;
  assign n12293 = n1746 & n7220;
  assign n12294 = x113 & n1750;
  assign n12295 = x112 & n1871;
  assign n12296 = ~n12294 & ~n12295;
  assign n12297 = x114 & n1873;
  assign n12298 = n12296 & ~n12297;
  assign n12299 = ~n12293 & n12298;
  assign n12300 = n12299 ^ x23;
  assign n12475 = n12474 ^ n12300;
  assign n12290 = n12197 ^ n12029;
  assign n12291 = ~n12198 & ~n12290;
  assign n12292 = n12291 ^ n12029;
  assign n12476 = n12475 ^ n12292;
  assign n12282 = n1404 & n7987;
  assign n12283 = x116 & n1408;
  assign n12284 = x115 & n1514;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = x117 & n1517;
  assign n12287 = n12285 & ~n12286;
  assign n12288 = ~n12282 & n12287;
  assign n12289 = n12288 ^ x20;
  assign n12477 = n12476 ^ n12289;
  assign n12279 = n12199 ^ n12018;
  assign n12280 = n12200 & n12279;
  assign n12281 = n12280 ^ n12018;
  assign n12478 = n12477 ^ n12281;
  assign n12271 = n1098 & n8820;
  assign n12272 = x119 & n1102;
  assign n12273 = x118 & n1198;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = x120 & n1201;
  assign n12276 = n12274 & ~n12275;
  assign n12277 = ~n12271 & n12276;
  assign n12278 = n12277 ^ x17;
  assign n12479 = n12478 ^ n12278;
  assign n12268 = n12201 ^ n12007;
  assign n12269 = ~n12202 & ~n12268;
  assign n12270 = n12269 ^ n12007;
  assign n12480 = n12479 ^ n12270;
  assign n12260 = n821 & n9691;
  assign n12261 = x121 & n898;
  assign n12262 = x123 & n901;
  assign n12263 = ~n12261 & ~n12262;
  assign n12264 = x122 & n824;
  assign n12265 = n12263 & ~n12264;
  assign n12266 = ~n12260 & n12265;
  assign n12267 = n12266 ^ x14;
  assign n12481 = n12480 ^ n12267;
  assign n12257 = n12203 ^ n11996;
  assign n12258 = n12204 & n12257;
  assign n12259 = n12258 ^ n11996;
  assign n12482 = n12481 ^ n12259;
  assign n12249 = n596 & ~n10570;
  assign n12250 = x124 & n673;
  assign n12251 = x126 & n676;
  assign n12252 = ~n12250 & ~n12251;
  assign n12253 = x125 & n601;
  assign n12254 = n12252 & ~n12253;
  assign n12255 = ~n12249 & n12254;
  assign n12256 = n12255 ^ x11;
  assign n12483 = n12482 ^ n12256;
  assign n12246 = n11993 ^ n11985;
  assign n12247 = n12206 & n12246;
  assign n12248 = n12247 ^ n12205;
  assign n12484 = n12483 ^ n12248;
  assign n12234 = n10278 ^ x8;
  assign n12235 = n12234 ^ x8;
  assign n12236 = ~x7 & x127;
  assign n12237 = n12236 ^ x8;
  assign n12238 = ~n12235 & ~n12237;
  assign n12239 = n12238 ^ x8;
  assign n12240 = ~n329 & ~n12239;
  assign n12241 = n340 ^ x7;
  assign n12242 = n398 & n12241;
  assign n12243 = x127 & n12242;
  assign n12244 = n12243 ^ x8;
  assign n12245 = ~n12240 & n12244;
  assign n12485 = n12484 ^ n12245;
  assign n12231 = n12207 ^ n11974;
  assign n12232 = n12208 & n12231;
  assign n12233 = n12232 ^ n11974;
  assign n12486 = n12485 ^ n12233;
  assign n12228 = n12209 ^ n11965;
  assign n12229 = ~n12210 & ~n12228;
  assign n12230 = n12229 ^ n11965;
  assign n12487 = n12486 ^ n12230;
  assign n12225 = n12223 ^ n11962;
  assign n12226 = ~n12212 & ~n12225;
  assign n12227 = n12226 ^ n12223;
  assign n12488 = n12487 ^ n12227;
  assign n12741 = n3585 & n4643;
  assign n12742 = x95 & n4653;
  assign n12743 = x96 & n4646;
  assign n12744 = ~n12742 & ~n12743;
  assign n12745 = x97 & n5046;
  assign n12746 = n12744 & ~n12745;
  assign n12747 = ~n12741 & n12746;
  assign n12748 = n12747 ^ x41;
  assign n12729 = n2607 & n5942;
  assign n12730 = x89 & n6186;
  assign n12731 = x90 & n5947;
  assign n12732 = ~n12730 & ~n12731;
  assign n12733 = x91 & n6406;
  assign n12734 = n12732 & ~n12733;
  assign n12735 = ~n12729 & n12734;
  assign n12736 = n12735 ^ x47;
  assign n12719 = n2176 & n6626;
  assign n12720 = x86 & n6884;
  assign n12721 = x88 & n6888;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = x87 & n6630;
  assign n12724 = n12722 & ~n12723;
  assign n12725 = ~n12719 & n12724;
  assign n12726 = n12725 ^ x50;
  assign n12705 = n1149 & n9002;
  assign n12706 = x77 & n9012;
  assign n12707 = x78 & n9005;
  assign n12708 = ~n12706 & ~n12707;
  assign n12709 = x79 & n9557;
  assign n12710 = n12708 & ~n12709;
  assign n12711 = ~n12705 & n12710;
  assign n12712 = n12711 ^ x59;
  assign n12702 = n12399 ^ n12391;
  assign n12703 = n12408 & n12702;
  assign n12704 = n12703 ^ n12407;
  assign n12713 = n12712 ^ n12704;
  assign n12680 = n12124 ^ x72;
  assign n12681 = n12680 ^ n12124;
  assign n12682 = n12124 ^ n10177;
  assign n12683 = n12682 ^ n12124;
  assign n12684 = ~n12681 & n12683;
  assign n12685 = n12684 ^ n12124;
  assign n12686 = x71 & n12685;
  assign n12687 = n12686 ^ n12124;
  assign n12688 = n12390 & ~n12687;
  assign n12689 = n10177 ^ x71;
  assign n12690 = n12379 ^ x72;
  assign n12691 = n12690 ^ n12689;
  assign n12692 = x70 ^ x63;
  assign n12693 = ~x70 & ~n12692;
  assign n12694 = n12693 ^ x72;
  assign n12695 = n12694 ^ x70;
  assign n12696 = n12691 & ~n12695;
  assign n12697 = n12696 ^ n12693;
  assign n12698 = n12697 ^ x70;
  assign n12699 = n12689 & ~n12698;
  assign n12700 = ~n12688 & ~n12699;
  assign n12671 = n870 & n9878;
  assign n12672 = x74 & n9888;
  assign n12673 = x76 & n10501;
  assign n12674 = ~n12672 & ~n12673;
  assign n12675 = x75 & n9881;
  assign n12676 = n12674 & ~n12675;
  assign n12677 = ~n12671 & n12676;
  assign n12678 = n12677 ^ x62;
  assign n12661 = x73 ^ x72;
  assign n12662 = n12661 ^ x63;
  assign n12663 = n12662 ^ n12661;
  assign n12664 = n12661 ^ n12379;
  assign n12665 = n12664 ^ n12661;
  assign n12666 = n12663 & n12665;
  assign n12667 = n12666 ^ n12661;
  assign n12668 = ~n10177 & n12667;
  assign n12669 = n12668 ^ n12661;
  assign n12670 = n12669 ^ x8;
  assign n12679 = n12678 ^ n12670;
  assign n12701 = n12700 ^ n12679;
  assign n12714 = n12713 ^ n12701;
  assign n12653 = n1454 & n8171;
  assign n12654 = x80 & n8181;
  assign n12655 = x82 & n8732;
  assign n12656 = ~n12654 & ~n12655;
  assign n12657 = x81 & n8174;
  assign n12658 = n12656 & ~n12657;
  assign n12659 = ~n12653 & n12658;
  assign n12660 = n12659 ^ x56;
  assign n12715 = n12714 ^ n12660;
  assign n12650 = n12378 ^ n12370;
  assign n12651 = ~n12410 & n12650;
  assign n12652 = n12651 ^ n12409;
  assign n12716 = n12715 ^ n12652;
  assign n12642 = n1801 & n7395;
  assign n12643 = x83 & n7650;
  assign n12644 = x84 & n7400;
  assign n12645 = ~n12643 & ~n12644;
  assign n12646 = x85 & n7652;
  assign n12647 = n12645 & ~n12646;
  assign n12648 = ~n12642 & n12647;
  assign n12649 = n12648 ^ x53;
  assign n12717 = n12716 ^ n12649;
  assign n12639 = n12411 ^ n12367;
  assign n12640 = n12420 & ~n12639;
  assign n12641 = n12640 ^ n12419;
  assign n12718 = n12717 ^ n12641;
  assign n12727 = n12726 ^ n12718;
  assign n12636 = n12421 ^ n12364;
  assign n12637 = n12430 & ~n12636;
  assign n12638 = n12637 ^ n12429;
  assign n12728 = n12727 ^ n12638;
  assign n12737 = n12736 ^ n12728;
  assign n12633 = n12434 ^ n12431;
  assign n12634 = n12443 & ~n12633;
  assign n12635 = n12634 ^ n12442;
  assign n12738 = n12737 ^ n12635;
  assign n12630 = n12444 ^ n12361;
  assign n12631 = n12453 & ~n12630;
  assign n12632 = n12631 ^ n12452;
  assign n12739 = n12738 ^ n12632;
  assign n12622 = n3078 & n5262;
  assign n12623 = x92 & n5488;
  assign n12624 = x94 & n5491;
  assign n12625 = ~n12623 & ~n12624;
  assign n12626 = x93 & n5266;
  assign n12627 = n12625 & ~n12626;
  assign n12628 = ~n12622 & n12627;
  assign n12629 = n12628 ^ x44;
  assign n12740 = n12739 ^ n12629;
  assign n12749 = n12748 ^ n12740;
  assign n12619 = n12462 ^ n12358;
  assign n12620 = ~n12463 & ~n12619;
  assign n12621 = n12620 ^ n12358;
  assign n12750 = n12749 ^ n12621;
  assign n12611 = n4040 & n4141;
  assign n12612 = x98 & n4267;
  assign n12613 = x99 & n4044;
  assign n12614 = ~n12612 & ~n12613;
  assign n12615 = x100 & n4270;
  assign n12616 = n12614 & ~n12615;
  assign n12617 = ~n12611 & n12616;
  assign n12618 = n12617 ^ x38;
  assign n12751 = n12750 ^ n12618;
  assign n12608 = n12464 ^ n12347;
  assign n12609 = n12465 & n12608;
  assign n12610 = n12609 ^ n12347;
  assign n12752 = n12751 ^ n12610;
  assign n12600 = n3522 & n4718;
  assign n12601 = x101 & n3699;
  assign n12602 = x103 & n3701;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = x102 & n3526;
  assign n12605 = n12603 & ~n12604;
  assign n12606 = ~n12600 & n12605;
  assign n12607 = n12606 ^ x35;
  assign n12753 = n12752 ^ n12607;
  assign n12597 = n12466 ^ n12336;
  assign n12598 = ~n12467 & ~n12597;
  assign n12599 = n12598 ^ n12336;
  assign n12754 = n12753 ^ n12599;
  assign n12589 = n3009 & n5351;
  assign n12590 = x104 & n3181;
  assign n12591 = x105 & n3013;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = x106 & n3183;
  assign n12594 = n12592 & ~n12593;
  assign n12595 = ~n12589 & n12594;
  assign n12596 = n12595 ^ x32;
  assign n12755 = n12754 ^ n12596;
  assign n12586 = n12468 ^ n12325;
  assign n12587 = n12469 & n12586;
  assign n12588 = n12587 ^ n12325;
  assign n12756 = n12755 ^ n12588;
  assign n12578 = n2527 & n6026;
  assign n12579 = x107 & n2690;
  assign n12580 = x109 & n2693;
  assign n12581 = ~n12579 & ~n12580;
  assign n12582 = x108 & n2530;
  assign n12583 = n12581 & ~n12582;
  assign n12584 = ~n12578 & n12583;
  assign n12585 = n12584 ^ x29;
  assign n12757 = n12756 ^ n12585;
  assign n12575 = n12470 ^ n12314;
  assign n12576 = ~n12471 & ~n12575;
  assign n12577 = n12576 ^ n12314;
  assign n12758 = n12757 ^ n12577;
  assign n12567 = n2102 & n6728;
  assign n12568 = x110 & n2112;
  assign n12569 = x112 & n2381;
  assign n12570 = ~n12568 & ~n12569;
  assign n12571 = x111 & n2105;
  assign n12572 = n12570 & ~n12571;
  assign n12573 = ~n12567 & n12572;
  assign n12574 = n12573 ^ x26;
  assign n12759 = n12758 ^ n12574;
  assign n12564 = n12472 ^ n12303;
  assign n12565 = n12473 & n12564;
  assign n12566 = n12565 ^ n12303;
  assign n12760 = n12759 ^ n12566;
  assign n12556 = n1746 & n7481;
  assign n12557 = x113 & n1871;
  assign n12558 = x114 & n1750;
  assign n12559 = ~n12557 & ~n12558;
  assign n12560 = x115 & n1873;
  assign n12561 = n12559 & ~n12560;
  assign n12562 = ~n12556 & n12561;
  assign n12563 = n12562 ^ x23;
  assign n12761 = n12760 ^ n12563;
  assign n12553 = n12474 ^ n12292;
  assign n12554 = ~n12475 & ~n12553;
  assign n12555 = n12554 ^ n12292;
  assign n12762 = n12761 ^ n12555;
  assign n12545 = n1404 & n8265;
  assign n12546 = x117 & n1408;
  assign n12547 = x116 & n1514;
  assign n12548 = ~n12546 & ~n12547;
  assign n12549 = x118 & n1517;
  assign n12550 = n12548 & ~n12549;
  assign n12551 = ~n12545 & n12550;
  assign n12552 = n12551 ^ x20;
  assign n12763 = n12762 ^ n12552;
  assign n12542 = n12476 ^ n12281;
  assign n12543 = n12477 & n12542;
  assign n12544 = n12543 ^ n12281;
  assign n12764 = n12763 ^ n12544;
  assign n12534 = n1098 & n9094;
  assign n12535 = x120 & n1102;
  assign n12536 = x119 & n1198;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = x121 & n1201;
  assign n12539 = n12537 & ~n12538;
  assign n12540 = ~n12534 & n12539;
  assign n12541 = n12540 ^ x17;
  assign n12765 = n12764 ^ n12541;
  assign n12531 = n12478 ^ n12270;
  assign n12532 = ~n12479 & ~n12531;
  assign n12533 = n12532 ^ n12270;
  assign n12766 = n12765 ^ n12533;
  assign n12523 = n821 & n9999;
  assign n12524 = x122 & n898;
  assign n12525 = x124 & n901;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = x123 & n824;
  assign n12528 = n12526 & ~n12527;
  assign n12529 = ~n12523 & n12528;
  assign n12530 = n12529 ^ x14;
  assign n12767 = n12766 ^ n12530;
  assign n12520 = n12480 ^ n12259;
  assign n12521 = n12481 & n12520;
  assign n12522 = n12521 ^ n12259;
  assign n12768 = n12767 ^ n12522;
  assign n12512 = n596 & ~n10855;
  assign n12513 = x125 & n673;
  assign n12514 = x126 & n601;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = x127 & n676;
  assign n12517 = n12515 & ~n12516;
  assign n12518 = ~n12512 & n12517;
  assign n12519 = n12518 ^ x11;
  assign n12769 = n12768 ^ n12519;
  assign n12509 = n12482 ^ n12248;
  assign n12510 = ~n12483 & n12509;
  assign n12511 = n12510 ^ n12248;
  assign n12770 = n12769 ^ n12511;
  assign n12491 = n12245 & ~n12484;
  assign n12492 = n12233 & n12491;
  assign n12489 = ~n12245 & n12484;
  assign n12490 = ~n12233 & n12489;
  assign n12493 = n12492 ^ n12490;
  assign n12494 = ~n12230 & n12493;
  assign n12495 = n12494 ^ n12492;
  assign n12496 = n12484 ^ n12233;
  assign n12497 = n12485 & ~n12496;
  assign n12498 = n12497 ^ n12233;
  assign n12499 = n12230 & n12498;
  assign n12500 = ~n12492 & ~n12499;
  assign n12501 = n12500 ^ n12227;
  assign n12502 = n12501 ^ n12500;
  assign n12503 = n12230 & ~n12490;
  assign n12504 = ~n12498 & ~n12503;
  assign n12505 = n12504 ^ n12500;
  assign n12506 = n12502 & ~n12505;
  assign n12507 = n12506 ^ n12500;
  assign n12508 = ~n12495 & n12507;
  assign n12771 = n12770 ^ n12508;
  assign n13017 = ~n12492 & n12770;
  assign n13018 = ~n12490 & ~n13017;
  assign n13019 = ~n12230 & ~n13018;
  assign n13020 = ~n12498 & n12770;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = ~n12227 & n13021;
  assign n13023 = n12230 & n13018;
  assign n13024 = n12498 & ~n12770;
  assign n13025 = ~n13023 & ~n13024;
  assign n13026 = ~n13022 & n13025;
  assign n12988 = n4040 & n4323;
  assign n12989 = x99 & n4267;
  assign n12990 = x100 & n4044;
  assign n12991 = ~n12989 & ~n12990;
  assign n12992 = x101 & n4270;
  assign n12993 = n12991 & ~n12992;
  assign n12994 = ~n12988 & n12993;
  assign n12995 = n12994 ^ x38;
  assign n12978 = n3763 & n4643;
  assign n12979 = x96 & n4653;
  assign n12980 = x97 & n4646;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = x98 & n5046;
  assign n12983 = n12981 & ~n12982;
  assign n12984 = ~n12978 & n12983;
  assign n12985 = n12984 ^ x41;
  assign n12968 = n3247 & n5262;
  assign n12969 = x93 & n5488;
  assign n12970 = x94 & n5266;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = x95 & n5491;
  assign n12973 = n12971 & ~n12972;
  assign n12974 = ~n12968 & n12973;
  assign n12975 = n12974 ^ x44;
  assign n12958 = n2755 & n5942;
  assign n12959 = x90 & n6186;
  assign n12960 = x91 & n5947;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = x92 & n6406;
  assign n12963 = n12961 & ~n12962;
  assign n12964 = ~n12958 & n12963;
  assign n12965 = n12964 ^ x47;
  assign n12948 = n2310 & n6626;
  assign n12949 = x88 & n6630;
  assign n12950 = x87 & n6884;
  assign n12951 = ~n12949 & ~n12950;
  assign n12952 = x89 & n6888;
  assign n12953 = n12951 & ~n12952;
  assign n12954 = ~n12948 & n12953;
  assign n12955 = n12954 ^ x50;
  assign n12938 = n1920 & n7395;
  assign n12939 = x85 & n7400;
  assign n12940 = x84 & n7650;
  assign n12941 = ~n12939 & ~n12940;
  assign n12942 = x86 & n7652;
  assign n12943 = n12941 & ~n12942;
  assign n12944 = ~n12938 & n12943;
  assign n12945 = n12944 ^ x53;
  assign n12935 = n12660 ^ n12652;
  assign n12936 = ~n12715 & n12935;
  assign n12937 = n12936 ^ n12714;
  assign n12946 = n12945 ^ n12937;
  assign n12925 = n1560 & n8171;
  assign n12926 = x81 & n8181;
  assign n12927 = x83 & n8732;
  assign n12928 = ~n12926 & ~n12927;
  assign n12929 = x82 & n8174;
  assign n12930 = n12928 & ~n12929;
  assign n12931 = ~n12925 & n12930;
  assign n12932 = n12931 ^ x56;
  assign n12915 = n1242 & n9002;
  assign n12916 = x78 & n9012;
  assign n12917 = x79 & n9005;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = x80 & n9557;
  assign n12920 = n12918 & ~n12919;
  assign n12921 = ~n12915 & n12920;
  assign n12922 = n12921 ^ x59;
  assign n12906 = n956 & n9878;
  assign n12907 = x75 & n9888;
  assign n12908 = x76 & n9881;
  assign n12909 = ~n12907 & ~n12908;
  assign n12910 = x77 & n10501;
  assign n12911 = n12909 & ~n12910;
  assign n12912 = ~n12906 & n12911;
  assign n12913 = n12912 ^ x62;
  assign n12902 = x74 & n10177;
  assign n12903 = x73 & n12123;
  assign n12904 = ~n12902 & ~n12903;
  assign n12893 = ~x62 & ~x63;
  assign n12894 = x72 ^ x8;
  assign n12895 = x73 ^ x71;
  assign n12896 = ~n12123 & n12895;
  assign n12897 = n12896 ^ x71;
  assign n12898 = n12897 ^ x72;
  assign n12899 = ~n12894 & n12898;
  assign n12900 = n12899 ^ x72;
  assign n12901 = ~n12893 & n12900;
  assign n12905 = n12904 ^ n12901;
  assign n12914 = n12913 ^ n12905;
  assign n12923 = n12922 ^ n12914;
  assign n12890 = n12700 ^ n12678;
  assign n12891 = ~n12679 & ~n12890;
  assign n12892 = n12891 ^ n12700;
  assign n12924 = n12923 ^ n12892;
  assign n12933 = n12932 ^ n12924;
  assign n12887 = n12712 ^ n12701;
  assign n12888 = n12713 & n12887;
  assign n12889 = n12888 ^ n12704;
  assign n12934 = n12933 ^ n12889;
  assign n12947 = n12946 ^ n12934;
  assign n12956 = n12955 ^ n12947;
  assign n12884 = n12716 ^ n12641;
  assign n12885 = ~n12717 & n12884;
  assign n12886 = n12885 ^ n12641;
  assign n12957 = n12956 ^ n12886;
  assign n12966 = n12965 ^ n12957;
  assign n12881 = n12726 ^ n12638;
  assign n12882 = ~n12727 & n12881;
  assign n12883 = n12882 ^ n12638;
  assign n12967 = n12966 ^ n12883;
  assign n12976 = n12975 ^ n12967;
  assign n12878 = n12736 ^ n12635;
  assign n12879 = ~n12737 & n12878;
  assign n12880 = n12879 ^ n12635;
  assign n12977 = n12976 ^ n12880;
  assign n12986 = n12985 ^ n12977;
  assign n12875 = n12738 ^ n12629;
  assign n12876 = n12739 & ~n12875;
  assign n12877 = n12876 ^ n12632;
  assign n12987 = n12986 ^ n12877;
  assign n12996 = n12995 ^ n12987;
  assign n12872 = n12748 ^ n12621;
  assign n12873 = ~n12749 & ~n12872;
  assign n12874 = n12873 ^ n12621;
  assign n12997 = n12996 ^ n12874;
  assign n12864 = n3522 & n4912;
  assign n12865 = x102 & n3699;
  assign n12866 = x103 & n3526;
  assign n12867 = ~n12865 & ~n12866;
  assign n12868 = x104 & n3701;
  assign n12869 = n12867 & ~n12868;
  assign n12870 = ~n12864 & n12869;
  assign n12871 = n12870 ^ x35;
  assign n12998 = n12997 ^ n12871;
  assign n12861 = n12750 ^ n12610;
  assign n12862 = n12751 & n12861;
  assign n12863 = n12862 ^ n12610;
  assign n12999 = n12998 ^ n12863;
  assign n12853 = n3009 & n5578;
  assign n12854 = x106 & n3013;
  assign n12855 = x105 & n3181;
  assign n12856 = ~n12854 & ~n12855;
  assign n12857 = x107 & n3183;
  assign n12858 = n12856 & ~n12857;
  assign n12859 = ~n12853 & n12858;
  assign n12860 = n12859 ^ x32;
  assign n13000 = n12999 ^ n12860;
  assign n12850 = n12752 ^ n12599;
  assign n12851 = ~n12753 & ~n12850;
  assign n12852 = n12851 ^ n12599;
  assign n13001 = n13000 ^ n12852;
  assign n12842 = n2527 & n6250;
  assign n12843 = x109 & n2530;
  assign n12844 = x108 & n2690;
  assign n12845 = ~n12843 & ~n12844;
  assign n12846 = x110 & n2693;
  assign n12847 = n12845 & ~n12846;
  assign n12848 = ~n12842 & n12847;
  assign n12849 = n12848 ^ x29;
  assign n13002 = n13001 ^ n12849;
  assign n12839 = n12754 ^ n12588;
  assign n12840 = n12755 & n12839;
  assign n12841 = n12840 ^ n12588;
  assign n13003 = n13002 ^ n12841;
  assign n12831 = n2102 & n6975;
  assign n12832 = x111 & n2112;
  assign n12833 = x113 & n2381;
  assign n12834 = ~n12832 & ~n12833;
  assign n12835 = x112 & n2105;
  assign n12836 = n12834 & ~n12835;
  assign n12837 = ~n12831 & n12836;
  assign n12838 = n12837 ^ x26;
  assign n13004 = n13003 ^ n12838;
  assign n12828 = n12756 ^ n12577;
  assign n12829 = ~n12757 & ~n12828;
  assign n12830 = n12829 ^ n12577;
  assign n13005 = n13004 ^ n12830;
  assign n12820 = n1746 & n7730;
  assign n12821 = x114 & n1871;
  assign n12822 = x115 & n1750;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = x116 & n1873;
  assign n12825 = n12823 & ~n12824;
  assign n12826 = ~n12820 & n12825;
  assign n12827 = n12826 ^ x23;
  assign n13006 = n13005 ^ n12827;
  assign n12817 = n12758 ^ n12566;
  assign n12818 = n12759 & n12817;
  assign n12819 = n12818 ^ n12566;
  assign n13007 = n13006 ^ n12819;
  assign n12809 = n1404 & n8542;
  assign n12810 = x117 & n1514;
  assign n12811 = x118 & n1408;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = x119 & n1517;
  assign n12814 = n12812 & ~n12813;
  assign n12815 = ~n12809 & n12814;
  assign n12816 = n12815 ^ x20;
  assign n13008 = n13007 ^ n12816;
  assign n12806 = n12760 ^ n12555;
  assign n12807 = ~n12761 & ~n12806;
  assign n12808 = n12807 ^ n12555;
  assign n13009 = n13008 ^ n12808;
  assign n12798 = n1098 & n9387;
  assign n12799 = x120 & n1198;
  assign n12800 = x121 & n1102;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = x122 & n1201;
  assign n12803 = n12801 & ~n12802;
  assign n12804 = ~n12798 & n12803;
  assign n12805 = n12804 ^ x17;
  assign n13010 = n13009 ^ n12805;
  assign n12795 = n12762 ^ n12544;
  assign n12796 = n12763 & n12795;
  assign n12797 = n12796 ^ n12544;
  assign n13011 = n13010 ^ n12797;
  assign n12787 = n821 & n10303;
  assign n12788 = x123 & n898;
  assign n12789 = x124 & n824;
  assign n12790 = ~n12788 & ~n12789;
  assign n12791 = x125 & n901;
  assign n12792 = n12790 & ~n12791;
  assign n12793 = ~n12787 & n12792;
  assign n12794 = n12793 ^ x14;
  assign n13012 = n13011 ^ n12794;
  assign n12784 = n12764 ^ n12533;
  assign n12785 = ~n12765 & ~n12784;
  assign n12786 = n12785 ^ n12533;
  assign n13013 = n13012 ^ n12786;
  assign n12778 = n596 & ~n10281;
  assign n12779 = x127 & n601;
  assign n12780 = x126 & n673;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = ~n12778 & n12781;
  assign n12783 = n12782 ^ x11;
  assign n13014 = n13013 ^ n12783;
  assign n12775 = n12766 ^ n12522;
  assign n12776 = n12767 & n12775;
  assign n12777 = n12776 ^ n12522;
  assign n13015 = n13014 ^ n12777;
  assign n12772 = n12519 ^ n12511;
  assign n12773 = n12769 & ~n12772;
  assign n12774 = n12773 ^ n12768;
  assign n13016 = n13015 ^ n12774;
  assign n13027 = n13026 ^ n13016;
  assign n13254 = n3522 & n5117;
  assign n13255 = x103 & n3699;
  assign n13256 = x104 & n3526;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = x105 & n3701;
  assign n13259 = n13257 & ~n13258;
  assign n13260 = ~n13254 & n13259;
  assign n13261 = n13260 ^ x35;
  assign n13245 = n4040 & n4509;
  assign n13246 = x100 & n4267;
  assign n13247 = x101 & n4044;
  assign n13248 = ~n13246 & ~n13247;
  assign n13249 = x102 & n4270;
  assign n13250 = n13248 & ~n13249;
  assign n13251 = ~n13245 & n13250;
  assign n13252 = n13251 ^ x38;
  assign n13235 = n3943 & n4643;
  assign n13236 = x97 & n4653;
  assign n13237 = x98 & n4646;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = x99 & n5046;
  assign n13240 = n13238 & ~n13239;
  assign n13241 = ~n13235 & n13240;
  assign n13242 = n13241 ^ x41;
  assign n13224 = n3403 & n5262;
  assign n13225 = x94 & n5488;
  assign n13226 = x96 & n5491;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = x95 & n5266;
  assign n13229 = n13227 & ~n13228;
  assign n13230 = ~n13224 & n13229;
  assign n13231 = n13230 ^ x44;
  assign n13214 = n2901 & n5942;
  assign n13215 = x91 & n6186;
  assign n13216 = x93 & n6406;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = x92 & n5947;
  assign n13219 = n13217 & ~n13218;
  assign n13220 = ~n13214 & n13219;
  assign n13221 = n13220 ^ x47;
  assign n13204 = n2448 & n6626;
  assign n13205 = x88 & n6884;
  assign n13206 = x89 & n6630;
  assign n13207 = ~n13205 & ~n13206;
  assign n13208 = x90 & n6888;
  assign n13209 = n13207 & ~n13208;
  assign n13210 = ~n13204 & n13209;
  assign n13211 = n13210 ^ x50;
  assign n13201 = n12945 ^ n12934;
  assign n13202 = ~n12946 & n13201;
  assign n13203 = n13202 ^ n12937;
  assign n13212 = n13211 ^ n13203;
  assign n13191 = n2039 & n7395;
  assign n13192 = x85 & n7650;
  assign n13193 = x87 & n7652;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = x86 & n7400;
  assign n13196 = n13194 & ~n13195;
  assign n13197 = ~n13191 & n13196;
  assign n13198 = n13197 ^ x53;
  assign n13181 = n1667 & n8171;
  assign n13182 = x82 & n8181;
  assign n13183 = x84 & n8732;
  assign n13184 = ~n13182 & ~n13183;
  assign n13185 = x83 & n8174;
  assign n13186 = n13184 & ~n13185;
  assign n13187 = ~n13181 & n13186;
  assign n13188 = n13187 ^ x56;
  assign n13166 = ~x75 & n12902;
  assign n13168 = x74 ^ x73;
  assign n13167 = ~x74 & x75;
  assign n13169 = n13168 ^ n13167;
  assign n13170 = n13169 ^ n13167;
  assign n13171 = n13167 ^ x63;
  assign n13172 = n13171 ^ n13167;
  assign n13173 = n13170 & n13172;
  assign n13174 = n13173 ^ n13167;
  assign n13175 = ~n10177 & n13174;
  assign n13176 = n13175 ^ n13167;
  assign n13177 = ~n13166 & ~n13176;
  assign n13163 = n12913 ^ n12901;
  assign n13164 = ~n12905 & ~n13163;
  assign n13165 = n13164 ^ n12913;
  assign n13178 = n13177 ^ n13165;
  assign n13155 = n1041 & n9878;
  assign n13156 = x76 & n9888;
  assign n13157 = x77 & n9881;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = x78 & n10501;
  assign n13160 = n13158 & ~n13159;
  assign n13161 = ~n13155 & n13160;
  assign n13162 = n13161 ^ x62;
  assign n13179 = n13178 ^ n13162;
  assign n13147 = n1340 & n9002;
  assign n13148 = x79 & n9012;
  assign n13149 = x80 & n9005;
  assign n13150 = ~n13148 & ~n13149;
  assign n13151 = x81 & n9557;
  assign n13152 = n13150 & ~n13151;
  assign n13153 = ~n13147 & n13152;
  assign n13154 = n13153 ^ x59;
  assign n13180 = n13179 ^ n13154;
  assign n13189 = n13188 ^ n13180;
  assign n13144 = n12922 ^ n12892;
  assign n13145 = ~n12923 & ~n13144;
  assign n13146 = n13145 ^ n12892;
  assign n13190 = n13189 ^ n13146;
  assign n13199 = n13198 ^ n13190;
  assign n13141 = n12932 ^ n12889;
  assign n13142 = n12933 & n13141;
  assign n13143 = n13142 ^ n12889;
  assign n13200 = n13199 ^ n13143;
  assign n13213 = n13212 ^ n13200;
  assign n13222 = n13221 ^ n13213;
  assign n13138 = n12947 ^ n12886;
  assign n13139 = n12956 & ~n13138;
  assign n13140 = n13139 ^ n12955;
  assign n13223 = n13222 ^ n13140;
  assign n13232 = n13231 ^ n13223;
  assign n13135 = n12957 ^ n12883;
  assign n13136 = n12966 & ~n13135;
  assign n13137 = n13136 ^ n12965;
  assign n13233 = n13232 ^ n13137;
  assign n13132 = n12967 ^ n12880;
  assign n13133 = n12976 & ~n13132;
  assign n13134 = n13133 ^ n12975;
  assign n13234 = n13233 ^ n13134;
  assign n13243 = n13242 ^ n13234;
  assign n13129 = n12977 ^ n12877;
  assign n13130 = n12986 & ~n13129;
  assign n13131 = n13130 ^ n12985;
  assign n13244 = n13243 ^ n13131;
  assign n13253 = n13252 ^ n13244;
  assign n13262 = n13261 ^ n13253;
  assign n13126 = n12995 ^ n12874;
  assign n13127 = ~n12996 & ~n13126;
  assign n13128 = n13127 ^ n12874;
  assign n13263 = n13262 ^ n13128;
  assign n13118 = n3009 & n5792;
  assign n13119 = x106 & n3181;
  assign n13120 = x107 & n3013;
  assign n13121 = ~n13119 & ~n13120;
  assign n13122 = x108 & n3183;
  assign n13123 = n13121 & ~n13122;
  assign n13124 = ~n13118 & n13123;
  assign n13125 = n13124 ^ x32;
  assign n13264 = n13263 ^ n13125;
  assign n13115 = n12997 ^ n12863;
  assign n13116 = n12998 & n13115;
  assign n13117 = n13116 ^ n12863;
  assign n13265 = n13264 ^ n13117;
  assign n13107 = n2527 & n6478;
  assign n13108 = x110 & n2530;
  assign n13109 = x109 & n2690;
  assign n13110 = ~n13108 & ~n13109;
  assign n13111 = x111 & n2693;
  assign n13112 = n13110 & ~n13111;
  assign n13113 = ~n13107 & n13112;
  assign n13114 = n13113 ^ x29;
  assign n13266 = n13265 ^ n13114;
  assign n13104 = n12999 ^ n12852;
  assign n13105 = ~n13000 & ~n13104;
  assign n13106 = n13105 ^ n12852;
  assign n13267 = n13266 ^ n13106;
  assign n13096 = n2102 & n7220;
  assign n13097 = x112 & n2112;
  assign n13098 = x113 & n2105;
  assign n13099 = ~n13097 & ~n13098;
  assign n13100 = x114 & n2381;
  assign n13101 = n13099 & ~n13100;
  assign n13102 = ~n13096 & n13101;
  assign n13103 = n13102 ^ x26;
  assign n13268 = n13267 ^ n13103;
  assign n13093 = n13001 ^ n12841;
  assign n13094 = n13002 & n13093;
  assign n13095 = n13094 ^ n12841;
  assign n13269 = n13268 ^ n13095;
  assign n13085 = n1746 & n7987;
  assign n13086 = x115 & n1871;
  assign n13087 = x116 & n1750;
  assign n13088 = ~n13086 & ~n13087;
  assign n13089 = x117 & n1873;
  assign n13090 = n13088 & ~n13089;
  assign n13091 = ~n13085 & n13090;
  assign n13092 = n13091 ^ x23;
  assign n13270 = n13269 ^ n13092;
  assign n13082 = n13003 ^ n12830;
  assign n13083 = ~n13004 & ~n13082;
  assign n13084 = n13083 ^ n12830;
  assign n13271 = n13270 ^ n13084;
  assign n13074 = n1404 & n8820;
  assign n13075 = x119 & n1408;
  assign n13076 = x118 & n1514;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = x120 & n1517;
  assign n13079 = n13077 & ~n13078;
  assign n13080 = ~n13074 & n13079;
  assign n13081 = n13080 ^ x20;
  assign n13272 = n13271 ^ n13081;
  assign n13071 = n13005 ^ n12819;
  assign n13072 = n13006 & n13071;
  assign n13073 = n13072 ^ n12819;
  assign n13273 = n13272 ^ n13073;
  assign n13063 = n1098 & n9691;
  assign n13064 = x122 & n1102;
  assign n13065 = x121 & n1198;
  assign n13066 = ~n13064 & ~n13065;
  assign n13067 = x123 & n1201;
  assign n13068 = n13066 & ~n13067;
  assign n13069 = ~n13063 & n13068;
  assign n13070 = n13069 ^ x17;
  assign n13274 = n13273 ^ n13070;
  assign n13060 = n13007 ^ n12808;
  assign n13061 = ~n13008 & ~n13060;
  assign n13062 = n13061 ^ n12808;
  assign n13275 = n13274 ^ n13062;
  assign n13052 = n821 & ~n10570;
  assign n13053 = x124 & n898;
  assign n13054 = x126 & n901;
  assign n13055 = ~n13053 & ~n13054;
  assign n13056 = x125 & n824;
  assign n13057 = n13055 & ~n13056;
  assign n13058 = ~n13052 & n13057;
  assign n13059 = n13058 ^ x14;
  assign n13276 = n13275 ^ n13059;
  assign n13049 = n13009 ^ n12797;
  assign n13050 = n13010 & n13049;
  assign n13051 = n13050 ^ n12797;
  assign n13277 = n13276 ^ n13051;
  assign n13037 = n10278 ^ x11;
  assign n13038 = n13037 ^ x11;
  assign n13039 = ~x10 & x127;
  assign n13040 = n13039 ^ x11;
  assign n13041 = ~n13038 & ~n13040;
  assign n13042 = n13041 ^ x11;
  assign n13043 = ~n534 & ~n13042;
  assign n13044 = n598 ^ x10;
  assign n13045 = n595 & n13044;
  assign n13046 = x127 & n13045;
  assign n13047 = n13046 ^ x11;
  assign n13048 = ~n13043 & n13047;
  assign n13278 = n13277 ^ n13048;
  assign n13034 = n13011 ^ n12786;
  assign n13035 = ~n13012 & ~n13034;
  assign n13036 = n13035 ^ n12786;
  assign n13279 = n13278 ^ n13036;
  assign n13031 = n13013 ^ n12777;
  assign n13032 = n13014 & n13031;
  assign n13033 = n13032 ^ n12777;
  assign n13280 = n13279 ^ n13033;
  assign n13028 = n13026 ^ n12774;
  assign n13029 = ~n13016 & n13028;
  assign n13030 = n13029 ^ n13026;
  assign n13281 = n13280 ^ n13030;
  assign n13496 = n3522 & n5351;
  assign n13497 = x104 & n3699;
  assign n13498 = x106 & n3701;
  assign n13499 = ~n13497 & ~n13498;
  assign n13500 = x105 & n3526;
  assign n13501 = n13499 & ~n13500;
  assign n13502 = ~n13496 & n13501;
  assign n13503 = n13502 ^ x35;
  assign n13484 = n4141 & n4643;
  assign n13485 = x98 & n4653;
  assign n13486 = x100 & n5046;
  assign n13487 = ~n13485 & ~n13486;
  assign n13488 = x99 & n4646;
  assign n13489 = n13487 & ~n13488;
  assign n13490 = ~n13484 & n13489;
  assign n13491 = n13490 ^ x41;
  assign n13474 = n3585 & n5262;
  assign n13475 = x95 & n5488;
  assign n13476 = x96 & n5266;
  assign n13477 = ~n13475 & ~n13476;
  assign n13478 = x97 & n5491;
  assign n13479 = n13477 & ~n13478;
  assign n13480 = ~n13474 & n13479;
  assign n13481 = n13480 ^ x44;
  assign n13464 = n3078 & n5942;
  assign n13465 = x92 & n6186;
  assign n13466 = x93 & n5947;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = x94 & n6406;
  assign n13469 = n13467 & ~n13468;
  assign n13470 = ~n13464 & n13469;
  assign n13471 = n13470 ^ x47;
  assign n13461 = n13213 ^ n13140;
  assign n13462 = n13222 & ~n13461;
  assign n13463 = n13462 ^ n13221;
  assign n13472 = n13471 ^ n13463;
  assign n13451 = n2607 & n6626;
  assign n13452 = x89 & n6884;
  assign n13453 = x90 & n6630;
  assign n13454 = ~n13452 & ~n13453;
  assign n13455 = x91 & n6888;
  assign n13456 = n13454 & ~n13455;
  assign n13457 = ~n13451 & n13456;
  assign n13458 = n13457 ^ x50;
  assign n13441 = n2176 & n7395;
  assign n13442 = x86 & n7650;
  assign n13443 = x87 & n7400;
  assign n13444 = ~n13442 & ~n13443;
  assign n13445 = x88 & n7652;
  assign n13446 = n13444 & ~n13445;
  assign n13447 = ~n13441 & n13446;
  assign n13448 = n13447 ^ x53;
  assign n13432 = n13165 & ~n13176;
  assign n13433 = ~x74 & n12903;
  assign n13434 = ~n13166 & ~n13433;
  assign n13435 = ~n13432 & n13434;
  assign n13423 = n1149 & n9878;
  assign n13424 = x77 & n9888;
  assign n13425 = x78 & n9881;
  assign n13426 = ~n13424 & ~n13425;
  assign n13427 = x79 & n10501;
  assign n13428 = n13426 & ~n13427;
  assign n13429 = ~n13423 & n13428;
  assign n13430 = n13429 ^ x62;
  assign n13413 = x76 ^ x63;
  assign n13414 = n13413 ^ x76;
  assign n13415 = x76 ^ x75;
  assign n13416 = n13415 ^ x76;
  assign n13417 = n13414 & n13416;
  assign n13418 = n13417 ^ x76;
  assign n13419 = ~n10177 & n13418;
  assign n13420 = n13419 ^ x76;
  assign n13421 = n13420 ^ n12904;
  assign n13422 = n13421 ^ x11;
  assign n13431 = n13430 ^ n13422;
  assign n13436 = n13435 ^ n13431;
  assign n13405 = n1454 & n9002;
  assign n13406 = x80 & n9012;
  assign n13407 = x81 & n9005;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = x82 & n9557;
  assign n13410 = n13408 & ~n13409;
  assign n13411 = ~n13405 & n13410;
  assign n13412 = n13411 ^ x59;
  assign n13437 = n13436 ^ n13412;
  assign n13402 = n13162 ^ n13154;
  assign n13403 = n13179 & ~n13402;
  assign n13404 = n13403 ^ n13178;
  assign n13438 = n13437 ^ n13404;
  assign n13394 = n1801 & n8171;
  assign n13395 = x83 & n8181;
  assign n13396 = x85 & n8732;
  assign n13397 = ~n13395 & ~n13396;
  assign n13398 = x84 & n8174;
  assign n13399 = n13397 & ~n13398;
  assign n13400 = ~n13394 & n13399;
  assign n13401 = n13400 ^ x56;
  assign n13439 = n13438 ^ n13401;
  assign n13391 = n13180 ^ n13146;
  assign n13392 = n13189 & n13391;
  assign n13393 = n13392 ^ n13188;
  assign n13440 = n13439 ^ n13393;
  assign n13449 = n13448 ^ n13440;
  assign n13388 = n13190 ^ n13143;
  assign n13389 = ~n13199 & n13388;
  assign n13390 = n13389 ^ n13198;
  assign n13450 = n13449 ^ n13390;
  assign n13459 = n13458 ^ n13450;
  assign n13385 = n13203 ^ n13200;
  assign n13386 = ~n13212 & ~n13385;
  assign n13387 = n13386 ^ n13211;
  assign n13460 = n13459 ^ n13387;
  assign n13473 = n13472 ^ n13460;
  assign n13482 = n13481 ^ n13473;
  assign n13382 = n13223 ^ n13137;
  assign n13383 = n13232 & ~n13382;
  assign n13384 = n13383 ^ n13231;
  assign n13483 = n13482 ^ n13384;
  assign n13492 = n13491 ^ n13483;
  assign n13379 = n13242 ^ n13233;
  assign n13380 = ~n13234 & n13379;
  assign n13381 = n13380 ^ n13242;
  assign n13493 = n13492 ^ n13381;
  assign n13376 = n13252 ^ n13131;
  assign n13377 = ~n13244 & n13376;
  assign n13378 = n13377 ^ n13252;
  assign n13494 = n13493 ^ n13378;
  assign n13368 = n4040 & n4718;
  assign n13369 = x101 & n4267;
  assign n13370 = x103 & n4270;
  assign n13371 = ~n13369 & ~n13370;
  assign n13372 = x102 & n4044;
  assign n13373 = n13371 & ~n13372;
  assign n13374 = ~n13368 & n13373;
  assign n13375 = n13374 ^ x38;
  assign n13495 = n13494 ^ n13375;
  assign n13504 = n13503 ^ n13495;
  assign n13365 = n13261 ^ n13128;
  assign n13366 = ~n13262 & ~n13365;
  assign n13367 = n13366 ^ n13128;
  assign n13505 = n13504 ^ n13367;
  assign n13357 = n3009 & n6026;
  assign n13358 = x108 & n3013;
  assign n13359 = x107 & n3181;
  assign n13360 = ~n13358 & ~n13359;
  assign n13361 = x109 & n3183;
  assign n13362 = n13360 & ~n13361;
  assign n13363 = ~n13357 & n13362;
  assign n13364 = n13363 ^ x32;
  assign n13506 = n13505 ^ n13364;
  assign n13354 = n13263 ^ n13117;
  assign n13355 = n13264 & n13354;
  assign n13356 = n13355 ^ n13117;
  assign n13507 = n13506 ^ n13356;
  assign n13346 = n2527 & n6728;
  assign n13347 = x110 & n2690;
  assign n13348 = x112 & n2693;
  assign n13349 = ~n13347 & ~n13348;
  assign n13350 = x111 & n2530;
  assign n13351 = n13349 & ~n13350;
  assign n13352 = ~n13346 & n13351;
  assign n13353 = n13352 ^ x29;
  assign n13508 = n13507 ^ n13353;
  assign n13343 = n13265 ^ n13106;
  assign n13344 = ~n13266 & ~n13343;
  assign n13345 = n13344 ^ n13106;
  assign n13509 = n13508 ^ n13345;
  assign n13335 = n2102 & n7481;
  assign n13336 = x113 & n2112;
  assign n13337 = x114 & n2105;
  assign n13338 = ~n13336 & ~n13337;
  assign n13339 = x115 & n2381;
  assign n13340 = n13338 & ~n13339;
  assign n13341 = ~n13335 & n13340;
  assign n13342 = n13341 ^ x26;
  assign n13510 = n13509 ^ n13342;
  assign n13332 = n13267 ^ n13095;
  assign n13333 = n13268 & n13332;
  assign n13334 = n13333 ^ n13095;
  assign n13511 = n13510 ^ n13334;
  assign n13324 = n1746 & n8265;
  assign n13325 = x116 & n1871;
  assign n13326 = x117 & n1750;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = x118 & n1873;
  assign n13329 = n13327 & ~n13328;
  assign n13330 = ~n13324 & n13329;
  assign n13331 = n13330 ^ x23;
  assign n13512 = n13511 ^ n13331;
  assign n13321 = n13269 ^ n13084;
  assign n13322 = ~n13270 & ~n13321;
  assign n13323 = n13322 ^ n13084;
  assign n13513 = n13512 ^ n13323;
  assign n13313 = n1404 & n9094;
  assign n13314 = x119 & n1514;
  assign n13315 = x121 & n1517;
  assign n13316 = ~n13314 & ~n13315;
  assign n13317 = x120 & n1408;
  assign n13318 = n13316 & ~n13317;
  assign n13319 = ~n13313 & n13318;
  assign n13320 = n13319 ^ x20;
  assign n13514 = n13513 ^ n13320;
  assign n13310 = n13271 ^ n13073;
  assign n13311 = n13272 & n13310;
  assign n13312 = n13311 ^ n13073;
  assign n13515 = n13514 ^ n13312;
  assign n13302 = n1098 & n9999;
  assign n13303 = x122 & n1198;
  assign n13304 = x123 & n1102;
  assign n13305 = ~n13303 & ~n13304;
  assign n13306 = x124 & n1201;
  assign n13307 = n13305 & ~n13306;
  assign n13308 = ~n13302 & n13307;
  assign n13309 = n13308 ^ x17;
  assign n13516 = n13515 ^ n13309;
  assign n13299 = n13273 ^ n13062;
  assign n13300 = ~n13274 & ~n13299;
  assign n13301 = n13300 ^ n13062;
  assign n13517 = n13516 ^ n13301;
  assign n13291 = n821 & ~n10855;
  assign n13292 = x125 & n898;
  assign n13293 = x126 & n824;
  assign n13294 = ~n13292 & ~n13293;
  assign n13295 = x127 & n901;
  assign n13296 = n13294 & ~n13295;
  assign n13297 = ~n13291 & n13296;
  assign n13298 = n13297 ^ x14;
  assign n13518 = n13517 ^ n13298;
  assign n13288 = n13275 ^ n13051;
  assign n13289 = n13276 & n13288;
  assign n13290 = n13289 ^ n13051;
  assign n13519 = n13518 ^ n13290;
  assign n13285 = n13277 ^ n13036;
  assign n13286 = n13278 & ~n13285;
  assign n13287 = n13286 ^ n13036;
  assign n13520 = n13519 ^ n13287;
  assign n13282 = n13033 ^ n13030;
  assign n13283 = n13280 & ~n13282;
  assign n13284 = n13283 ^ n13030;
  assign n13521 = n13520 ^ n13284;
  assign n13733 = n3009 & n6250;
  assign n13734 = x108 & n3181;
  assign n13735 = x109 & n3013;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = x110 & n3183;
  assign n13738 = n13736 & ~n13737;
  assign n13739 = ~n13733 & n13738;
  assign n13740 = n13739 ^ x32;
  assign n13724 = n3522 & n5578;
  assign n13725 = x105 & n3699;
  assign n13726 = x106 & n3526;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = x107 & n3701;
  assign n13729 = n13727 & ~n13728;
  assign n13730 = ~n13724 & n13729;
  assign n13731 = n13730 ^ x35;
  assign n13714 = n4040 & n4912;
  assign n13715 = x102 & n4267;
  assign n13716 = x104 & n4270;
  assign n13717 = ~n13715 & ~n13716;
  assign n13718 = x103 & n4044;
  assign n13719 = n13717 & ~n13718;
  assign n13720 = ~n13714 & n13719;
  assign n13721 = n13720 ^ x38;
  assign n13704 = n4323 & n4643;
  assign n13705 = x99 & n4653;
  assign n13706 = x100 & n4646;
  assign n13707 = ~n13705 & ~n13706;
  assign n13708 = x101 & n5046;
  assign n13709 = n13707 & ~n13708;
  assign n13710 = ~n13704 & n13709;
  assign n13711 = n13710 ^ x41;
  assign n13693 = n3763 & n5262;
  assign n13694 = x96 & n5488;
  assign n13695 = x98 & n5491;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = x97 & n5266;
  assign n13698 = n13696 & ~n13697;
  assign n13699 = ~n13693 & n13698;
  assign n13700 = n13699 ^ x44;
  assign n13683 = n3247 & n5942;
  assign n13684 = x93 & n6186;
  assign n13685 = x95 & n6406;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = x94 & n5947;
  assign n13688 = n13686 & ~n13687;
  assign n13689 = ~n13683 & n13688;
  assign n13690 = n13689 ^ x47;
  assign n13673 = n2755 & n6626;
  assign n13674 = x90 & n6884;
  assign n13675 = x92 & n6888;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = x91 & n6630;
  assign n13678 = n13676 & ~n13677;
  assign n13679 = ~n13673 & n13678;
  assign n13680 = n13679 ^ x50;
  assign n13663 = n2310 & n7395;
  assign n13664 = x88 & n7400;
  assign n13665 = x87 & n7650;
  assign n13666 = ~n13664 & ~n13665;
  assign n13667 = x89 & n7652;
  assign n13668 = n13666 & ~n13667;
  assign n13669 = ~n13663 & n13668;
  assign n13670 = n13669 ^ x53;
  assign n13653 = n1920 & n8171;
  assign n13654 = x85 & n8174;
  assign n13655 = x84 & n8181;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = x86 & n8732;
  assign n13658 = n13656 & ~n13657;
  assign n13659 = ~n13653 & n13658;
  assign n13660 = n13659 ^ x56;
  assign n13650 = n13436 ^ n13404;
  assign n13651 = ~n13437 & n13650;
  assign n13652 = n13651 ^ n13404;
  assign n13661 = n13660 ^ n13652;
  assign n13640 = n1560 & n9002;
  assign n13641 = x81 & n9012;
  assign n13642 = x83 & n9557;
  assign n13643 = ~n13641 & ~n13642;
  assign n13644 = x82 & n9005;
  assign n13645 = n13643 & ~n13644;
  assign n13646 = ~n13640 & n13645;
  assign n13647 = n13646 ^ x59;
  assign n13631 = n1242 & n9878;
  assign n13632 = x78 & n9888;
  assign n13633 = x80 & n10501;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = x79 & n9881;
  assign n13636 = n13634 & ~n13635;
  assign n13637 = ~n13631 & n13636;
  assign n13638 = n13637 ^ x62;
  assign n13622 = x77 ^ x63;
  assign n13623 = n13622 ^ x77;
  assign n13624 = x77 ^ x76;
  assign n13625 = n13624 ^ x77;
  assign n13626 = n13623 & n13625;
  assign n13627 = n13626 ^ x77;
  assign n13628 = ~n10177 & n13627;
  assign n13629 = n13628 ^ x77;
  assign n13619 = n12904 ^ x11;
  assign n13620 = n13421 & n13619;
  assign n13621 = n13620 ^ x11;
  assign n13630 = n13629 ^ n13621;
  assign n13639 = n13638 ^ n13630;
  assign n13648 = n13647 ^ n13639;
  assign n13616 = n13435 ^ n13430;
  assign n13617 = n13431 & ~n13616;
  assign n13618 = n13617 ^ n13435;
  assign n13649 = n13648 ^ n13618;
  assign n13662 = n13661 ^ n13649;
  assign n13671 = n13670 ^ n13662;
  assign n13613 = n13438 ^ n13393;
  assign n13614 = ~n13439 & n13613;
  assign n13615 = n13614 ^ n13393;
  assign n13672 = n13671 ^ n13615;
  assign n13681 = n13680 ^ n13672;
  assign n13610 = n13448 ^ n13390;
  assign n13611 = ~n13449 & n13610;
  assign n13612 = n13611 ^ n13390;
  assign n13682 = n13681 ^ n13612;
  assign n13691 = n13690 ^ n13682;
  assign n13607 = n13458 ^ n13387;
  assign n13608 = ~n13459 & n13607;
  assign n13609 = n13608 ^ n13387;
  assign n13692 = n13691 ^ n13609;
  assign n13701 = n13700 ^ n13692;
  assign n13604 = n13471 ^ n13460;
  assign n13605 = n13472 & ~n13604;
  assign n13606 = n13605 ^ n13463;
  assign n13702 = n13701 ^ n13606;
  assign n13601 = n13481 ^ n13384;
  assign n13602 = ~n13482 & n13601;
  assign n13603 = n13602 ^ n13384;
  assign n13703 = n13702 ^ n13603;
  assign n13712 = n13711 ^ n13703;
  assign n13598 = n13491 ^ n13381;
  assign n13599 = ~n13492 & n13598;
  assign n13600 = n13599 ^ n13381;
  assign n13713 = n13712 ^ n13600;
  assign n13722 = n13721 ^ n13713;
  assign n13595 = n13493 ^ n13375;
  assign n13596 = n13494 & ~n13595;
  assign n13597 = n13596 ^ n13378;
  assign n13723 = n13722 ^ n13597;
  assign n13732 = n13731 ^ n13723;
  assign n13741 = n13740 ^ n13732;
  assign n13592 = n13503 ^ n13367;
  assign n13593 = ~n13504 & ~n13592;
  assign n13594 = n13593 ^ n13367;
  assign n13742 = n13741 ^ n13594;
  assign n13589 = n13505 ^ n13356;
  assign n13590 = n13506 & n13589;
  assign n13591 = n13590 ^ n13356;
  assign n13743 = n13742 ^ n13591;
  assign n13581 = n2527 & n6975;
  assign n13582 = x111 & n2690;
  assign n13583 = x113 & n2693;
  assign n13584 = ~n13582 & ~n13583;
  assign n13585 = x112 & n2530;
  assign n13586 = n13584 & ~n13585;
  assign n13587 = ~n13581 & n13586;
  assign n13588 = n13587 ^ x29;
  assign n13744 = n13743 ^ n13588;
  assign n13573 = n2102 & n7730;
  assign n13574 = x114 & n2112;
  assign n13575 = x116 & n2381;
  assign n13576 = ~n13574 & ~n13575;
  assign n13577 = x115 & n2105;
  assign n13578 = n13576 & ~n13577;
  assign n13579 = ~n13573 & n13578;
  assign n13580 = n13579 ^ x26;
  assign n13745 = n13744 ^ n13580;
  assign n13570 = n13507 ^ n13345;
  assign n13571 = ~n13508 & ~n13570;
  assign n13572 = n13571 ^ n13345;
  assign n13746 = n13745 ^ n13572;
  assign n13562 = n1746 & n8542;
  assign n13563 = x117 & n1871;
  assign n13564 = x119 & n1873;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = x118 & n1750;
  assign n13567 = n13565 & ~n13566;
  assign n13568 = ~n13562 & n13567;
  assign n13569 = n13568 ^ x23;
  assign n13747 = n13746 ^ n13569;
  assign n13559 = n13509 ^ n13334;
  assign n13560 = n13510 & n13559;
  assign n13561 = n13560 ^ n13334;
  assign n13748 = n13747 ^ n13561;
  assign n13551 = n1404 & n9387;
  assign n13552 = x121 & n1408;
  assign n13553 = x120 & n1514;
  assign n13554 = ~n13552 & ~n13553;
  assign n13555 = x122 & n1517;
  assign n13556 = n13554 & ~n13555;
  assign n13557 = ~n13551 & n13556;
  assign n13558 = n13557 ^ x20;
  assign n13749 = n13748 ^ n13558;
  assign n13548 = n13511 ^ n13323;
  assign n13549 = ~n13512 & ~n13548;
  assign n13550 = n13549 ^ n13323;
  assign n13750 = n13749 ^ n13550;
  assign n13540 = n1098 & n10303;
  assign n13541 = x124 & n1102;
  assign n13542 = x123 & n1198;
  assign n13543 = ~n13541 & ~n13542;
  assign n13544 = x125 & n1201;
  assign n13545 = n13543 & ~n13544;
  assign n13546 = ~n13540 & n13545;
  assign n13547 = n13546 ^ x17;
  assign n13751 = n13750 ^ n13547;
  assign n13537 = n13513 ^ n13312;
  assign n13538 = n13514 & n13537;
  assign n13539 = n13538 ^ n13312;
  assign n13752 = n13751 ^ n13539;
  assign n13531 = n821 & ~n10281;
  assign n13532 = x126 & n898;
  assign n13533 = x127 & n824;
  assign n13534 = ~n13532 & ~n13533;
  assign n13535 = ~n13531 & n13534;
  assign n13536 = n13535 ^ x14;
  assign n13753 = n13752 ^ n13536;
  assign n13528 = n13515 ^ n13301;
  assign n13529 = ~n13516 & ~n13528;
  assign n13530 = n13529 ^ n13301;
  assign n13754 = n13753 ^ n13530;
  assign n13525 = n13517 ^ n13290;
  assign n13526 = n13518 & n13525;
  assign n13527 = n13526 ^ n13290;
  assign n13755 = n13754 ^ n13527;
  assign n13522 = n13287 ^ n13284;
  assign n13523 = n13520 & ~n13522;
  assign n13524 = n13523 ^ n13284;
  assign n13756 = n13755 ^ n13524;
  assign n13975 = n3009 & n6478;
  assign n13976 = x109 & n3181;
  assign n13977 = x110 & n3013;
  assign n13978 = ~n13976 & ~n13977;
  assign n13979 = x111 & n3183;
  assign n13980 = n13978 & ~n13979;
  assign n13981 = ~n13975 & n13980;
  assign n13982 = n13981 ^ x32;
  assign n13965 = n3522 & n5792;
  assign n13966 = x106 & n3699;
  assign n13967 = x107 & n3526;
  assign n13968 = ~n13966 & ~n13967;
  assign n13969 = x108 & n3701;
  assign n13970 = n13968 & ~n13969;
  assign n13971 = ~n13965 & n13970;
  assign n13972 = n13971 ^ x35;
  assign n13955 = n4040 & n5117;
  assign n13956 = x103 & n4267;
  assign n13957 = x105 & n4270;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = x104 & n4044;
  assign n13960 = n13958 & ~n13959;
  assign n13961 = ~n13955 & n13960;
  assign n13962 = n13961 ^ x38;
  assign n13945 = n4509 & n4643;
  assign n13946 = x100 & n4653;
  assign n13947 = x102 & n5046;
  assign n13948 = ~n13946 & ~n13947;
  assign n13949 = x101 & n4646;
  assign n13950 = n13948 & ~n13949;
  assign n13951 = ~n13945 & n13950;
  assign n13952 = n13951 ^ x41;
  assign n13934 = n3943 & n5262;
  assign n13935 = x97 & n5488;
  assign n13936 = x98 & n5266;
  assign n13937 = ~n13935 & ~n13936;
  assign n13938 = x99 & n5491;
  assign n13939 = n13937 & ~n13938;
  assign n13940 = ~n13934 & n13939;
  assign n13941 = n13940 ^ x44;
  assign n13924 = n3403 & n5942;
  assign n13925 = x94 & n6186;
  assign n13926 = x96 & n6406;
  assign n13927 = ~n13925 & ~n13926;
  assign n13928 = x95 & n5947;
  assign n13929 = n13927 & ~n13928;
  assign n13930 = ~n13924 & n13929;
  assign n13931 = n13930 ^ x47;
  assign n13914 = n2901 & n6626;
  assign n13915 = x91 & n6884;
  assign n13916 = x93 & n6888;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = x92 & n6630;
  assign n13919 = n13917 & ~n13918;
  assign n13920 = ~n13914 & n13919;
  assign n13921 = n13920 ^ x50;
  assign n13904 = n2448 & n7395;
  assign n13905 = x88 & n7650;
  assign n13906 = x89 & n7400;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = x90 & n7652;
  assign n13909 = n13907 & ~n13908;
  assign n13910 = ~n13904 & n13909;
  assign n13911 = n13910 ^ x53;
  assign n13901 = n13660 ^ n13649;
  assign n13902 = n13661 & n13901;
  assign n13903 = n13902 ^ n13652;
  assign n13912 = n13911 ^ n13903;
  assign n13891 = n2039 & n8171;
  assign n13892 = x85 & n8181;
  assign n13893 = x86 & n8174;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = x87 & n8732;
  assign n13896 = n13894 & ~n13895;
  assign n13897 = ~n13891 & n13896;
  assign n13898 = n13897 ^ x56;
  assign n13882 = n1667 & n9002;
  assign n13883 = x82 & n9012;
  assign n13884 = x84 & n9557;
  assign n13885 = ~n13883 & ~n13884;
  assign n13886 = x83 & n9005;
  assign n13887 = n13885 & ~n13886;
  assign n13888 = ~n13882 & n13887;
  assign n13889 = n13888 ^ x59;
  assign n13873 = n1340 & n9878;
  assign n13874 = x79 & n9888;
  assign n13875 = x81 & n10501;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = x80 & n9881;
  assign n13878 = n13876 & ~n13877;
  assign n13879 = ~n13873 & n13878;
  assign n13862 = n859 ^ x62;
  assign n13863 = n13862 ^ x63;
  assign n13864 = n13863 ^ n859;
  assign n13865 = n13624 ^ n859;
  assign n13866 = n13865 ^ n859;
  assign n13867 = n859 ^ x63;
  assign n13868 = n13867 ^ n859;
  assign n13869 = n13866 & n13868;
  assign n13870 = n13869 ^ n859;
  assign n13871 = ~n13864 & n13870;
  assign n13872 = n13871 ^ n13862;
  assign n13880 = n13879 ^ n13872;
  assign n13859 = n13638 ^ n13621;
  assign n13860 = ~n13630 & n13859;
  assign n13861 = n13860 ^ n13638;
  assign n13881 = n13880 ^ n13861;
  assign n13890 = n13889 ^ n13881;
  assign n13899 = n13898 ^ n13890;
  assign n13856 = n13647 ^ n13618;
  assign n13857 = ~n13648 & ~n13856;
  assign n13858 = n13857 ^ n13618;
  assign n13900 = n13899 ^ n13858;
  assign n13913 = n13912 ^ n13900;
  assign n13922 = n13921 ^ n13913;
  assign n13853 = n13662 ^ n13615;
  assign n13854 = ~n13671 & n13853;
  assign n13855 = n13854 ^ n13670;
  assign n13923 = n13922 ^ n13855;
  assign n13932 = n13931 ^ n13923;
  assign n13850 = n13672 ^ n13612;
  assign n13851 = ~n13681 & n13850;
  assign n13852 = n13851 ^ n13680;
  assign n13933 = n13932 ^ n13852;
  assign n13942 = n13941 ^ n13933;
  assign n13847 = n13682 ^ n13609;
  assign n13848 = ~n13691 & n13847;
  assign n13849 = n13848 ^ n13690;
  assign n13943 = n13942 ^ n13849;
  assign n13844 = n13692 ^ n13606;
  assign n13845 = ~n13701 & n13844;
  assign n13846 = n13845 ^ n13700;
  assign n13944 = n13943 ^ n13846;
  assign n13953 = n13952 ^ n13944;
  assign n13841 = n13711 ^ n13603;
  assign n13842 = n13703 & n13841;
  assign n13843 = n13842 ^ n13711;
  assign n13954 = n13953 ^ n13843;
  assign n13963 = n13962 ^ n13954;
  assign n13838 = n13721 ^ n13600;
  assign n13839 = n13713 & n13838;
  assign n13840 = n13839 ^ n13721;
  assign n13964 = n13963 ^ n13840;
  assign n13973 = n13972 ^ n13964;
  assign n13835 = n13731 ^ n13597;
  assign n13836 = n13723 & n13835;
  assign n13837 = n13836 ^ n13731;
  assign n13974 = n13973 ^ n13837;
  assign n13983 = n13982 ^ n13974;
  assign n13832 = n13740 ^ n13594;
  assign n13833 = n13741 & ~n13832;
  assign n13834 = n13833 ^ n13594;
  assign n13984 = n13983 ^ n13834;
  assign n13824 = n2527 & n7220;
  assign n13825 = x112 & n2690;
  assign n13826 = x114 & n2693;
  assign n13827 = ~n13825 & ~n13826;
  assign n13828 = x113 & n2530;
  assign n13829 = n13827 & ~n13828;
  assign n13830 = ~n13824 & n13829;
  assign n13831 = n13830 ^ x29;
  assign n13985 = n13984 ^ n13831;
  assign n13821 = n13742 ^ n13588;
  assign n13822 = ~n13743 & ~n13821;
  assign n13823 = n13822 ^ n13591;
  assign n13986 = n13985 ^ n13823;
  assign n13813 = n2102 & n7987;
  assign n13814 = x115 & n2112;
  assign n13815 = x116 & n2105;
  assign n13816 = ~n13814 & ~n13815;
  assign n13817 = x117 & n2381;
  assign n13818 = n13816 & ~n13817;
  assign n13819 = ~n13813 & n13818;
  assign n13820 = n13819 ^ x26;
  assign n13987 = n13986 ^ n13820;
  assign n13805 = n1746 & n8820;
  assign n13806 = x119 & n1750;
  assign n13807 = x118 & n1871;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = x120 & n1873;
  assign n13810 = n13808 & ~n13809;
  assign n13811 = ~n13805 & n13810;
  assign n13812 = n13811 ^ x23;
  assign n13988 = n13987 ^ n13812;
  assign n13802 = n13744 ^ n13572;
  assign n13803 = n13745 & n13802;
  assign n13804 = n13803 ^ n13572;
  assign n13989 = n13988 ^ n13804;
  assign n13799 = n13746 ^ n13561;
  assign n13800 = ~n13747 & ~n13799;
  assign n13801 = n13800 ^ n13561;
  assign n13990 = n13989 ^ n13801;
  assign n13791 = n1404 & n9691;
  assign n13792 = x121 & n1514;
  assign n13793 = x123 & n1517;
  assign n13794 = ~n13792 & ~n13793;
  assign n13795 = x122 & n1408;
  assign n13796 = n13794 & ~n13795;
  assign n13797 = ~n13791 & n13796;
  assign n13798 = n13797 ^ x20;
  assign n13991 = n13990 ^ n13798;
  assign n13788 = n13748 ^ n13550;
  assign n13789 = n13749 & n13788;
  assign n13790 = n13789 ^ n13550;
  assign n13992 = n13991 ^ n13790;
  assign n13780 = n1098 & ~n10570;
  assign n13781 = x125 & n1102;
  assign n13782 = x124 & n1198;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = x126 & n1201;
  assign n13785 = n13783 & ~n13784;
  assign n13786 = ~n13780 & n13785;
  assign n13787 = n13786 ^ x17;
  assign n13993 = n13992 ^ n13787;
  assign n13766 = x127 & n813;
  assign n13767 = ~x14 & ~n13766;
  assign n13768 = n13767 ^ x13;
  assign n13769 = n666 & n11409;
  assign n13770 = n13769 ^ n13767;
  assign n13771 = ~n13767 & n13770;
  assign n13772 = n13771 ^ n13767;
  assign n13773 = x127 & n897;
  assign n13774 = ~n13772 & ~n13773;
  assign n13775 = n13774 ^ n13771;
  assign n13776 = n13775 ^ n13767;
  assign n13777 = n13776 ^ n13769;
  assign n13778 = ~n13768 & n13777;
  assign n13779 = n13778 ^ x13;
  assign n13994 = n13993 ^ n13779;
  assign n13763 = n13750 ^ n13539;
  assign n13764 = ~n13751 & ~n13763;
  assign n13765 = n13764 ^ n13539;
  assign n13995 = n13994 ^ n13765;
  assign n13760 = n13752 ^ n13530;
  assign n13761 = n13753 & n13760;
  assign n13762 = n13761 ^ n13530;
  assign n13996 = n13995 ^ n13762;
  assign n13757 = n13527 ^ n13524;
  assign n13758 = n13755 & ~n13757;
  assign n13759 = n13758 ^ n13524;
  assign n13997 = n13996 ^ n13759;
  assign n14233 = n2102 & n8265;
  assign n14234 = x116 & n2112;
  assign n14235 = x117 & n2105;
  assign n14236 = ~n14234 & ~n14235;
  assign n14237 = x118 & n2381;
  assign n14238 = n14236 & ~n14237;
  assign n14239 = ~n14233 & n14238;
  assign n14240 = n14239 ^ x26;
  assign n14223 = n2527 & n7481;
  assign n14224 = x114 & n2530;
  assign n14225 = x113 & n2690;
  assign n14226 = ~n14224 & ~n14225;
  assign n14227 = x115 & n2693;
  assign n14228 = n14226 & ~n14227;
  assign n14229 = ~n14223 & n14228;
  assign n14230 = n14229 ^ x29;
  assign n14213 = n3009 & n6728;
  assign n14214 = x110 & n3181;
  assign n14215 = x111 & n3013;
  assign n14216 = ~n14214 & ~n14215;
  assign n14217 = x112 & n3183;
  assign n14218 = n14216 & ~n14217;
  assign n14219 = ~n14213 & n14218;
  assign n14220 = n14219 ^ x32;
  assign n14203 = n3522 & n6026;
  assign n14204 = x107 & n3699;
  assign n14205 = x109 & n3701;
  assign n14206 = ~n14204 & ~n14205;
  assign n14207 = x108 & n3526;
  assign n14208 = n14206 & ~n14207;
  assign n14209 = ~n14203 & n14208;
  assign n14210 = n14209 ^ x35;
  assign n14193 = n4040 & n5351;
  assign n14194 = x104 & n4267;
  assign n14195 = x106 & n4270;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = x105 & n4044;
  assign n14198 = n14196 & ~n14197;
  assign n14199 = ~n14193 & n14198;
  assign n14200 = n14199 ^ x38;
  assign n14183 = n4643 & n4718;
  assign n14184 = x101 & n4653;
  assign n14185 = x102 & n4646;
  assign n14186 = ~n14184 & ~n14185;
  assign n14187 = x103 & n5046;
  assign n14188 = n14186 & ~n14187;
  assign n14189 = ~n14183 & n14188;
  assign n14190 = n14189 ^ x41;
  assign n14173 = n4141 & n5262;
  assign n14174 = x98 & n5488;
  assign n14175 = x100 & n5491;
  assign n14176 = ~n14174 & ~n14175;
  assign n14177 = x99 & n5266;
  assign n14178 = n14176 & ~n14177;
  assign n14179 = ~n14173 & n14178;
  assign n14180 = n14179 ^ x44;
  assign n14163 = n3585 & n5942;
  assign n14164 = x95 & n6186;
  assign n14165 = x97 & n6406;
  assign n14166 = ~n14164 & ~n14165;
  assign n14167 = x96 & n5947;
  assign n14168 = n14166 & ~n14167;
  assign n14169 = ~n14163 & n14168;
  assign n14170 = n14169 ^ x47;
  assign n14153 = n3078 & n6626;
  assign n14154 = x92 & n6884;
  assign n14155 = x94 & n6888;
  assign n14156 = ~n14154 & ~n14155;
  assign n14157 = x93 & n6630;
  assign n14158 = n14156 & ~n14157;
  assign n14159 = ~n14153 & n14158;
  assign n14160 = n14159 ^ x50;
  assign n14143 = n2607 & n7395;
  assign n14144 = x90 & n7400;
  assign n14145 = x89 & n7650;
  assign n14146 = ~n14144 & ~n14145;
  assign n14147 = x91 & n7652;
  assign n14148 = n14146 & ~n14147;
  assign n14149 = ~n14143 & n14148;
  assign n14150 = n14149 ^ x53;
  assign n14133 = n2176 & n8171;
  assign n14134 = x86 & n8181;
  assign n14135 = x87 & n8174;
  assign n14136 = ~n14134 & ~n14135;
  assign n14137 = x88 & n8732;
  assign n14138 = n14136 & ~n14137;
  assign n14139 = ~n14133 & n14138;
  assign n14140 = n14139 ^ x56;
  assign n14123 = n1801 & n9002;
  assign n14124 = x83 & n9012;
  assign n14125 = x84 & n9005;
  assign n14126 = ~n14124 & ~n14125;
  assign n14127 = x85 & n9557;
  assign n14128 = n14126 & ~n14127;
  assign n14129 = ~n14123 & n14128;
  assign n14130 = n14129 ^ x59;
  assign n14105 = x63 & n859;
  assign n14106 = ~n13879 & ~n14105;
  assign n14107 = ~x77 & x78;
  assign n14108 = x63 & n14107;
  assign n14109 = ~x62 & ~n14108;
  assign n14110 = ~n14106 & n14109;
  assign n14111 = n13879 ^ x77;
  assign n14112 = ~n13624 & n14111;
  assign n14113 = n14112 ^ x77;
  assign n14114 = n12123 & ~n14113;
  assign n14115 = ~n14110 & ~n14114;
  assign n14116 = x62 & ~x63;
  assign n14117 = n13879 ^ x78;
  assign n14118 = ~n859 & n14117;
  assign n14119 = n14118 ^ x78;
  assign n14120 = n14116 & ~n14119;
  assign n14121 = n14115 & ~n14120;
  assign n14096 = n1454 & n9878;
  assign n14097 = x80 & n9888;
  assign n14098 = x81 & n9881;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = x82 & n10501;
  assign n14101 = n14099 & ~n14100;
  assign n14102 = ~n14096 & n14101;
  assign n14103 = n14102 ^ x62;
  assign n14087 = x79 ^ x63;
  assign n14088 = n14087 ^ x79;
  assign n14089 = n934 ^ x79;
  assign n14090 = n14088 & n14089;
  assign n14091 = n14090 ^ x79;
  assign n14092 = ~n10177 & n14091;
  assign n14093 = n14092 ^ x79;
  assign n14094 = n14093 ^ x14;
  assign n14095 = n14094 ^ n13629;
  assign n14104 = n14103 ^ n14095;
  assign n14122 = n14121 ^ n14104;
  assign n14131 = n14130 ^ n14122;
  assign n14084 = n13889 ^ n13861;
  assign n14085 = n13881 & n14084;
  assign n14086 = n14085 ^ n13889;
  assign n14132 = n14131 ^ n14086;
  assign n14141 = n14140 ^ n14132;
  assign n14081 = n13890 ^ n13858;
  assign n14082 = ~n13899 & ~n14081;
  assign n14083 = n14082 ^ n13898;
  assign n14142 = n14141 ^ n14083;
  assign n14151 = n14150 ^ n14142;
  assign n14078 = n13903 ^ n13900;
  assign n14079 = n13912 & ~n14078;
  assign n14080 = n14079 ^ n13911;
  assign n14152 = n14151 ^ n14080;
  assign n14161 = n14160 ^ n14152;
  assign n14075 = n13913 ^ n13855;
  assign n14076 = n13922 & ~n14075;
  assign n14077 = n14076 ^ n13921;
  assign n14162 = n14161 ^ n14077;
  assign n14171 = n14170 ^ n14162;
  assign n14072 = n13923 ^ n13852;
  assign n14073 = n13932 & ~n14072;
  assign n14074 = n14073 ^ n13931;
  assign n14172 = n14171 ^ n14074;
  assign n14181 = n14180 ^ n14172;
  assign n14069 = n13933 ^ n13849;
  assign n14070 = n13942 & ~n14069;
  assign n14071 = n14070 ^ n13941;
  assign n14182 = n14181 ^ n14071;
  assign n14191 = n14190 ^ n14182;
  assign n14066 = n13952 ^ n13943;
  assign n14067 = ~n13944 & n14066;
  assign n14068 = n14067 ^ n13952;
  assign n14192 = n14191 ^ n14068;
  assign n14201 = n14200 ^ n14192;
  assign n14063 = n13962 ^ n13953;
  assign n14064 = ~n13954 & n14063;
  assign n14065 = n14064 ^ n13962;
  assign n14202 = n14201 ^ n14065;
  assign n14211 = n14210 ^ n14202;
  assign n14060 = n13972 ^ n13963;
  assign n14061 = ~n13964 & n14060;
  assign n14062 = n14061 ^ n13972;
  assign n14212 = n14211 ^ n14062;
  assign n14221 = n14220 ^ n14212;
  assign n14057 = n13982 ^ n13837;
  assign n14058 = ~n13974 & n14057;
  assign n14059 = n14058 ^ n13982;
  assign n14222 = n14221 ^ n14059;
  assign n14231 = n14230 ^ n14222;
  assign n14054 = n13983 ^ n13831;
  assign n14055 = ~n13984 & ~n14054;
  assign n14056 = n14055 ^ n13834;
  assign n14232 = n14231 ^ n14056;
  assign n14241 = n14240 ^ n14232;
  assign n14051 = n13985 ^ n13820;
  assign n14052 = n13986 & n14051;
  assign n14053 = n14052 ^ n13823;
  assign n14242 = n14241 ^ n14053;
  assign n14043 = n1746 & n9094;
  assign n14044 = x119 & n1871;
  assign n14045 = x120 & n1750;
  assign n14046 = ~n14044 & ~n14045;
  assign n14047 = x121 & n1873;
  assign n14048 = n14046 & ~n14047;
  assign n14049 = ~n14043 & n14048;
  assign n14050 = n14049 ^ x23;
  assign n14243 = n14242 ^ n14050;
  assign n14040 = n13987 ^ n13804;
  assign n14041 = ~n13988 & ~n14040;
  assign n14042 = n14041 ^ n13804;
  assign n14244 = n14243 ^ n14042;
  assign n14032 = n1404 & n9999;
  assign n14033 = x123 & n1408;
  assign n14034 = x122 & n1514;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = x124 & n1517;
  assign n14037 = n14035 & ~n14036;
  assign n14038 = ~n14032 & n14037;
  assign n14039 = n14038 ^ x20;
  assign n14245 = n14244 ^ n14039;
  assign n14029 = n13989 ^ n13798;
  assign n14030 = n13990 & n14029;
  assign n14031 = n14030 ^ n13801;
  assign n14246 = n14245 ^ n14031;
  assign n14021 = n1098 & ~n10855;
  assign n14022 = x126 & n1102;
  assign n14023 = x125 & n1198;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = x127 & n1201;
  assign n14026 = n14024 & ~n14025;
  assign n14027 = ~n14021 & n14026;
  assign n14028 = n14027 ^ x17;
  assign n14247 = n14246 ^ n14028;
  assign n14018 = n13991 ^ n13787;
  assign n14019 = ~n13992 & ~n14018;
  assign n14020 = n14019 ^ n13790;
  assign n14248 = n14247 ^ n14020;
  assign n14000 = n13779 & n13993;
  assign n14001 = n13765 & n14000;
  assign n13998 = ~n13779 & ~n13993;
  assign n13999 = ~n13765 & n13998;
  assign n14002 = n14001 ^ n13999;
  assign n14003 = ~n13762 & n14002;
  assign n14004 = n14003 ^ n14001;
  assign n14005 = ~n13762 & ~n14001;
  assign n14006 = n13993 ^ n13765;
  assign n14007 = ~n13994 & n14006;
  assign n14008 = n14007 ^ n13765;
  assign n14009 = ~n14005 & n14008;
  assign n14010 = n14009 ^ n13759;
  assign n14011 = n14010 ^ n14009;
  assign n14012 = n13762 & ~n13999;
  assign n14013 = ~n14008 & ~n14012;
  assign n14014 = n14013 ^ n14009;
  assign n14015 = n14011 & n14014;
  assign n14016 = n14015 ^ n14009;
  assign n14017 = ~n14004 & ~n14016;
  assign n14249 = n14248 ^ n14017;
  assign n14466 = n13762 & n13765;
  assign n14467 = ~n13998 & n14466;
  assign n14468 = n14248 & ~n14467;
  assign n14469 = ~n13759 & ~n14468;
  assign n14470 = ~n13762 & ~n13765;
  assign n14471 = ~n14248 & ~n14470;
  assign n14472 = ~n14000 & ~n14471;
  assign n14473 = ~n14469 & n14472;
  assign n14474 = ~n13998 & ~n14248;
  assign n14475 = n13765 ^ n13762;
  assign n14476 = n13762 ^ n13759;
  assign n14477 = n14475 & ~n14476;
  assign n14478 = n14477 ^ n13762;
  assign n14479 = ~n14474 & ~n14478;
  assign n14480 = ~n14473 & ~n14479;
  assign n14449 = n2102 & n8542;
  assign n14450 = x117 & n2112;
  assign n14451 = x118 & n2105;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = x119 & n2381;
  assign n14454 = n14452 & ~n14453;
  assign n14455 = ~n14449 & n14454;
  assign n14456 = n14455 ^ x26;
  assign n14440 = n2527 & n7730;
  assign n14441 = x115 & n2530;
  assign n14442 = x114 & n2690;
  assign n14443 = ~n14441 & ~n14442;
  assign n14444 = x116 & n2693;
  assign n14445 = n14443 & ~n14444;
  assign n14446 = ~n14440 & n14445;
  assign n14447 = n14446 ^ x29;
  assign n14430 = n3009 & n6975;
  assign n14431 = x111 & n3181;
  assign n14432 = x112 & n3013;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = x113 & n3183;
  assign n14435 = n14433 & ~n14434;
  assign n14436 = ~n14430 & n14435;
  assign n14437 = n14436 ^ x32;
  assign n14419 = n3522 & n6250;
  assign n14420 = x108 & n3699;
  assign n14421 = x110 & n3701;
  assign n14422 = ~n14420 & ~n14421;
  assign n14423 = x109 & n3526;
  assign n14424 = n14422 & ~n14423;
  assign n14425 = ~n14419 & n14424;
  assign n14426 = n14425 ^ x35;
  assign n14416 = n14200 ^ n14065;
  assign n14417 = n14201 & n14416;
  assign n14418 = n14417 ^ n14065;
  assign n14427 = n14426 ^ n14418;
  assign n14407 = n4040 & n5578;
  assign n14408 = x105 & n4267;
  assign n14409 = x106 & n4044;
  assign n14410 = ~n14408 & ~n14409;
  assign n14411 = x107 & n4270;
  assign n14412 = n14410 & ~n14411;
  assign n14413 = ~n14407 & n14412;
  assign n14414 = n14413 ^ x38;
  assign n14397 = n4643 & n4912;
  assign n14398 = x102 & n4653;
  assign n14399 = x103 & n4646;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = x104 & n5046;
  assign n14402 = n14400 & ~n14401;
  assign n14403 = ~n14397 & n14402;
  assign n14404 = n14403 ^ x41;
  assign n14386 = n4323 & n5262;
  assign n14387 = x99 & n5488;
  assign n14388 = x101 & n5491;
  assign n14389 = ~n14387 & ~n14388;
  assign n14390 = x100 & n5266;
  assign n14391 = n14389 & ~n14390;
  assign n14392 = ~n14386 & n14391;
  assign n14393 = n14392 ^ x44;
  assign n14383 = n14170 ^ n14074;
  assign n14384 = n14171 & n14383;
  assign n14385 = n14384 ^ n14074;
  assign n14394 = n14393 ^ n14385;
  assign n14373 = n3763 & n5942;
  assign n14374 = x96 & n6186;
  assign n14375 = x98 & n6406;
  assign n14376 = ~n14374 & ~n14375;
  assign n14377 = x97 & n5947;
  assign n14378 = n14376 & ~n14377;
  assign n14379 = ~n14373 & n14378;
  assign n14380 = n14379 ^ x47;
  assign n14363 = n3247 & n6626;
  assign n14364 = x93 & n6884;
  assign n14365 = x94 & n6630;
  assign n14366 = ~n14364 & ~n14365;
  assign n14367 = x95 & n6888;
  assign n14368 = n14366 & ~n14367;
  assign n14369 = ~n14363 & n14368;
  assign n14370 = n14369 ^ x50;
  assign n14353 = n2755 & n7395;
  assign n14354 = x91 & n7400;
  assign n14355 = x90 & n7650;
  assign n14356 = ~n14354 & ~n14355;
  assign n14357 = x92 & n7652;
  assign n14358 = n14356 & ~n14357;
  assign n14359 = ~n14353 & n14358;
  assign n14360 = n14359 ^ x53;
  assign n14350 = n14140 ^ n14083;
  assign n14351 = n14141 & n14350;
  assign n14352 = n14351 ^ n14083;
  assign n14361 = n14360 ^ n14352;
  assign n14340 = n2310 & n8171;
  assign n14341 = x87 & n8181;
  assign n14342 = x89 & n8732;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = x88 & n8174;
  assign n14345 = n14343 & ~n14344;
  assign n14346 = ~n14340 & n14345;
  assign n14347 = n14346 ^ x56;
  assign n14337 = n14130 ^ n14086;
  assign n14338 = n14131 & n14337;
  assign n14339 = n14338 ^ n14086;
  assign n14348 = n14347 ^ n14339;
  assign n14327 = n1920 & n9002;
  assign n14328 = x84 & n9012;
  assign n14329 = x86 & n9557;
  assign n14330 = ~n14328 & ~n14329;
  assign n14331 = x85 & n9005;
  assign n14332 = n14330 & ~n14331;
  assign n14333 = ~n14327 & n14332;
  assign n14334 = n14333 ^ x59;
  assign n14319 = n1560 & n9878;
  assign n14320 = x81 & n9888;
  assign n14321 = x83 & n10501;
  assign n14322 = ~n14320 & ~n14321;
  assign n14323 = x82 & n9881;
  assign n14324 = n14322 & ~n14323;
  assign n14325 = ~n14319 & n14324;
  assign n14314 = n13629 ^ x14;
  assign n14315 = n14093 ^ n13629;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = n14316 ^ x14;
  assign n14310 = x63 & x80;
  assign n14308 = ~x63 & n1030;
  assign n14309 = n14308 ^ x79;
  assign n14311 = n14310 ^ n14309;
  assign n14312 = ~x62 & ~n14311;
  assign n14313 = n14312 ^ n14309;
  assign n14318 = n14317 ^ n14313;
  assign n14326 = n14325 ^ n14318;
  assign n14335 = n14334 ^ n14326;
  assign n14305 = n14121 ^ n14103;
  assign n14306 = ~n14104 & ~n14305;
  assign n14307 = n14306 ^ n14121;
  assign n14336 = n14335 ^ n14307;
  assign n14349 = n14348 ^ n14336;
  assign n14362 = n14361 ^ n14349;
  assign n14371 = n14370 ^ n14362;
  assign n14302 = n14150 ^ n14080;
  assign n14303 = n14151 & n14302;
  assign n14304 = n14303 ^ n14080;
  assign n14372 = n14371 ^ n14304;
  assign n14381 = n14380 ^ n14372;
  assign n14299 = n14160 ^ n14077;
  assign n14300 = n14161 & n14299;
  assign n14301 = n14300 ^ n14077;
  assign n14382 = n14381 ^ n14301;
  assign n14395 = n14394 ^ n14382;
  assign n14296 = n14180 ^ n14071;
  assign n14297 = n14181 & n14296;
  assign n14298 = n14297 ^ n14071;
  assign n14396 = n14395 ^ n14298;
  assign n14405 = n14404 ^ n14396;
  assign n14293 = n14182 ^ n14068;
  assign n14294 = ~n14191 & n14293;
  assign n14295 = n14294 ^ n14190;
  assign n14406 = n14405 ^ n14295;
  assign n14415 = n14414 ^ n14406;
  assign n14428 = n14427 ^ n14415;
  assign n14290 = n14210 ^ n14062;
  assign n14291 = n14211 & n14290;
  assign n14292 = n14291 ^ n14062;
  assign n14429 = n14428 ^ n14292;
  assign n14438 = n14437 ^ n14429;
  assign n14287 = n14220 ^ n14059;
  assign n14288 = n14221 & n14287;
  assign n14289 = n14288 ^ n14059;
  assign n14439 = n14438 ^ n14289;
  assign n14448 = n14447 ^ n14439;
  assign n14457 = n14456 ^ n14448;
  assign n14284 = n14230 ^ n14056;
  assign n14285 = n14231 & ~n14284;
  assign n14286 = n14285 ^ n14056;
  assign n14458 = n14457 ^ n14286;
  assign n14281 = n14240 ^ n14053;
  assign n14282 = ~n14241 & ~n14281;
  assign n14283 = n14282 ^ n14053;
  assign n14459 = n14458 ^ n14283;
  assign n14273 = n1746 & n9387;
  assign n14274 = x121 & n1750;
  assign n14275 = x120 & n1871;
  assign n14276 = ~n14274 & ~n14275;
  assign n14277 = x122 & n1873;
  assign n14278 = n14276 & ~n14277;
  assign n14279 = ~n14273 & n14278;
  assign n14280 = n14279 ^ x23;
  assign n14460 = n14459 ^ n14280;
  assign n14270 = n14242 ^ n14042;
  assign n14271 = n14243 & n14270;
  assign n14272 = n14271 ^ n14042;
  assign n14461 = n14460 ^ n14272;
  assign n14262 = n1404 & n10303;
  assign n14263 = x123 & n1514;
  assign n14264 = x124 & n1408;
  assign n14265 = ~n14263 & ~n14264;
  assign n14266 = x125 & n1517;
  assign n14267 = n14265 & ~n14266;
  assign n14268 = ~n14262 & n14267;
  assign n14269 = n14268 ^ x20;
  assign n14462 = n14461 ^ n14269;
  assign n14259 = n14244 ^ n14031;
  assign n14260 = ~n14245 & ~n14259;
  assign n14261 = n14260 ^ n14031;
  assign n14463 = n14462 ^ n14261;
  assign n14253 = n1098 & ~n10281;
  assign n14254 = x126 & n1198;
  assign n14255 = x127 & n1102;
  assign n14256 = ~n14254 & ~n14255;
  assign n14257 = ~n14253 & n14256;
  assign n14258 = n14257 ^ x17;
  assign n14464 = n14463 ^ n14258;
  assign n14250 = n14246 ^ n14020;
  assign n14251 = n14247 & n14250;
  assign n14252 = n14251 ^ n14020;
  assign n14465 = n14464 ^ n14252;
  assign n14481 = n14480 ^ n14465;
  assign n14709 = n14252 & n14261;
  assign n14710 = n14258 & ~n14462;
  assign n14716 = n14709 & ~n14710;
  assign n14712 = ~n14252 & ~n14261;
  assign n14713 = ~n14258 & n14462;
  assign n14717 = ~n14712 & n14713;
  assign n14718 = ~n14716 & ~n14717;
  assign n14711 = ~n14709 & n14710;
  assign n14714 = n14712 & ~n14713;
  assign n14715 = ~n14711 & ~n14714;
  assign n14719 = n14718 ^ n14715;
  assign n14720 = ~n14480 & n14719;
  assign n14721 = n14720 ^ n14718;
  assign n14722 = n14261 ^ n14252;
  assign n14723 = n14713 ^ n14710;
  assign n14724 = n14710 ^ n14261;
  assign n14725 = n14724 ^ n14710;
  assign n14726 = n14723 & n14725;
  assign n14727 = n14726 ^ n14710;
  assign n14728 = ~n14722 & n14727;
  assign n14729 = n14721 & ~n14728;
  assign n14698 = n1404 & ~n10570;
  assign n14699 = x124 & n1514;
  assign n14700 = x125 & n1408;
  assign n14701 = ~n14699 & ~n14700;
  assign n14702 = x126 & n1517;
  assign n14703 = n14701 & ~n14702;
  assign n14704 = ~n14698 & n14703;
  assign n14705 = n14704 ^ x20;
  assign n14688 = n1746 & n9691;
  assign n14689 = x122 & n1750;
  assign n14690 = x121 & n1871;
  assign n14691 = ~n14689 & ~n14690;
  assign n14692 = x123 & n1873;
  assign n14693 = n14691 & ~n14692;
  assign n14694 = ~n14688 & n14693;
  assign n14695 = n14694 ^ x23;
  assign n14678 = n2102 & n8820;
  assign n14679 = x118 & n2112;
  assign n14680 = x119 & n2105;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = x120 & n2381;
  assign n14683 = n14681 & ~n14682;
  assign n14684 = ~n14678 & n14683;
  assign n14685 = n14684 ^ x26;
  assign n14668 = n2527 & n7987;
  assign n14669 = x115 & n2690;
  assign n14670 = x116 & n2530;
  assign n14671 = ~n14669 & ~n14670;
  assign n14672 = x117 & n2693;
  assign n14673 = n14671 & ~n14672;
  assign n14674 = ~n14668 & n14673;
  assign n14675 = n14674 ^ x29;
  assign n14658 = n3009 & n7220;
  assign n14659 = x113 & n3013;
  assign n14660 = x112 & n3181;
  assign n14661 = ~n14659 & ~n14660;
  assign n14662 = x114 & n3183;
  assign n14663 = n14661 & ~n14662;
  assign n14664 = ~n14658 & n14663;
  assign n14665 = n14664 ^ x32;
  assign n14648 = n3522 & n6478;
  assign n14649 = x109 & n3699;
  assign n14650 = x111 & n3701;
  assign n14651 = ~n14649 & ~n14650;
  assign n14652 = x110 & n3526;
  assign n14653 = n14651 & ~n14652;
  assign n14654 = ~n14648 & n14653;
  assign n14655 = n14654 ^ x35;
  assign n14638 = n4040 & n5792;
  assign n14639 = x106 & n4267;
  assign n14640 = x108 & n4270;
  assign n14641 = ~n14639 & ~n14640;
  assign n14642 = x107 & n4044;
  assign n14643 = n14641 & ~n14642;
  assign n14644 = ~n14638 & n14643;
  assign n14645 = n14644 ^ x38;
  assign n14628 = n4643 & n5117;
  assign n14629 = x103 & n4653;
  assign n14630 = x104 & n4646;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = x105 & n5046;
  assign n14633 = n14631 & ~n14632;
  assign n14634 = ~n14628 & n14633;
  assign n14635 = n14634 ^ x41;
  assign n14617 = n4509 & n5262;
  assign n14618 = x100 & n5488;
  assign n14619 = x101 & n5266;
  assign n14620 = ~n14618 & ~n14619;
  assign n14621 = x102 & n5491;
  assign n14622 = n14620 & ~n14621;
  assign n14623 = ~n14617 & n14622;
  assign n14624 = n14623 ^ x44;
  assign n14607 = n3943 & n5942;
  assign n14608 = x97 & n6186;
  assign n14609 = x98 & n5947;
  assign n14610 = ~n14608 & ~n14609;
  assign n14611 = x99 & n6406;
  assign n14612 = n14610 & ~n14611;
  assign n14613 = ~n14607 & n14612;
  assign n14614 = n14613 ^ x47;
  assign n14604 = n14362 ^ n14304;
  assign n14605 = n14371 & ~n14604;
  assign n14606 = n14605 ^ n14370;
  assign n14615 = n14614 ^ n14606;
  assign n14594 = n3403 & n6626;
  assign n14595 = x94 & n6884;
  assign n14596 = x95 & n6630;
  assign n14597 = ~n14595 & ~n14596;
  assign n14598 = x96 & n6888;
  assign n14599 = n14597 & ~n14598;
  assign n14600 = ~n14594 & n14599;
  assign n14601 = n14600 ^ x50;
  assign n14584 = n2901 & n7395;
  assign n14585 = x91 & n7650;
  assign n14586 = x92 & n7400;
  assign n14587 = ~n14585 & ~n14586;
  assign n14588 = x93 & n7652;
  assign n14589 = n14587 & ~n14588;
  assign n14590 = ~n14584 & n14589;
  assign n14591 = n14590 ^ x53;
  assign n14575 = n2448 & n8171;
  assign n14576 = x88 & n8181;
  assign n14577 = x90 & n8732;
  assign n14578 = ~n14576 & ~n14577;
  assign n14579 = x89 & n8174;
  assign n14580 = n14578 & ~n14579;
  assign n14581 = ~n14575 & n14580;
  assign n14582 = n14581 ^ x56;
  assign n14565 = n2039 & n9002;
  assign n14566 = x85 & n9012;
  assign n14567 = x87 & n9557;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = x86 & n9005;
  assign n14570 = n14568 & ~n14569;
  assign n14571 = ~n14565 & n14570;
  assign n14572 = n14571 ^ x59;
  assign n14556 = n1667 & n9878;
  assign n14557 = x82 & n9888;
  assign n14558 = x84 & n10501;
  assign n14559 = ~n14557 & ~n14558;
  assign n14560 = x83 & n9881;
  assign n14561 = n14559 & ~n14560;
  assign n14562 = ~n14556 & n14561;
  assign n14545 = n1130 ^ x62;
  assign n14546 = n14545 ^ x63;
  assign n14547 = n14546 ^ n1130;
  assign n14548 = n1130 ^ x63;
  assign n14549 = n14548 ^ n1130;
  assign n14550 = n1130 ^ n1030;
  assign n14551 = n14550 ^ n1130;
  assign n14552 = n14549 & n14551;
  assign n14553 = n14552 ^ n1130;
  assign n14554 = ~n14547 & n14553;
  assign n14555 = n14554 ^ n14545;
  assign n14563 = n14562 ^ n14555;
  assign n14535 = n14325 ^ n14317;
  assign n14539 = n14325 ^ n14310;
  assign n14540 = n14535 & n14539;
  assign n14541 = n14540 ^ n14325;
  assign n14536 = n14325 ^ n14309;
  assign n14537 = ~n14535 & ~n14536;
  assign n14538 = n14537 ^ n14325;
  assign n14542 = n14541 ^ n14538;
  assign n14543 = x62 & ~n14542;
  assign n14544 = n14543 ^ n14541;
  assign n14564 = n14563 ^ n14544;
  assign n14573 = n14572 ^ n14564;
  assign n14532 = n14326 ^ n14307;
  assign n14533 = ~n14335 & ~n14532;
  assign n14534 = n14533 ^ n14334;
  assign n14574 = n14573 ^ n14534;
  assign n14583 = n14582 ^ n14574;
  assign n14592 = n14591 ^ n14583;
  assign n14529 = n14339 ^ n14336;
  assign n14530 = n14348 & ~n14529;
  assign n14531 = n14530 ^ n14347;
  assign n14593 = n14592 ^ n14531;
  assign n14602 = n14601 ^ n14593;
  assign n14526 = n14360 ^ n14349;
  assign n14527 = n14361 & ~n14526;
  assign n14528 = n14527 ^ n14352;
  assign n14603 = n14602 ^ n14528;
  assign n14616 = n14615 ^ n14603;
  assign n14625 = n14624 ^ n14616;
  assign n14523 = n14372 ^ n14301;
  assign n14524 = n14381 & ~n14523;
  assign n14525 = n14524 ^ n14380;
  assign n14626 = n14625 ^ n14525;
  assign n14520 = n14385 ^ n14382;
  assign n14521 = n14394 & ~n14520;
  assign n14522 = n14521 ^ n14393;
  assign n14627 = n14626 ^ n14522;
  assign n14636 = n14635 ^ n14627;
  assign n14517 = n14404 ^ n14298;
  assign n14518 = ~n14396 & n14517;
  assign n14519 = n14518 ^ n14404;
  assign n14637 = n14636 ^ n14519;
  assign n14646 = n14645 ^ n14637;
  assign n14514 = n14414 ^ n14295;
  assign n14515 = ~n14406 & n14514;
  assign n14516 = n14515 ^ n14414;
  assign n14647 = n14646 ^ n14516;
  assign n14656 = n14655 ^ n14647;
  assign n14511 = n14426 ^ n14415;
  assign n14512 = n14427 & ~n14511;
  assign n14513 = n14512 ^ n14418;
  assign n14657 = n14656 ^ n14513;
  assign n14666 = n14665 ^ n14657;
  assign n14508 = n14437 ^ n14428;
  assign n14509 = ~n14429 & n14508;
  assign n14510 = n14509 ^ n14437;
  assign n14667 = n14666 ^ n14510;
  assign n14676 = n14675 ^ n14667;
  assign n14505 = n14447 ^ n14289;
  assign n14506 = ~n14439 & n14505;
  assign n14507 = n14506 ^ n14447;
  assign n14677 = n14676 ^ n14507;
  assign n14686 = n14685 ^ n14677;
  assign n14502 = n14456 ^ n14286;
  assign n14503 = ~n14457 & ~n14502;
  assign n14504 = n14503 ^ n14286;
  assign n14687 = n14686 ^ n14504;
  assign n14696 = n14695 ^ n14687;
  assign n14499 = n14458 ^ n14280;
  assign n14500 = n14459 & n14499;
  assign n14501 = n14500 ^ n14283;
  assign n14697 = n14696 ^ n14501;
  assign n14706 = n14705 ^ n14697;
  assign n14485 = x127 & n1001;
  assign n14486 = ~x17 & ~n14485;
  assign n14487 = n14486 ^ x16;
  assign n14488 = n907 & n11409;
  assign n14489 = n14488 ^ n14486;
  assign n14490 = ~n14486 & n14489;
  assign n14491 = n14490 ^ n14486;
  assign n14492 = x127 & n1197;
  assign n14493 = ~n14491 & ~n14492;
  assign n14494 = n14493 ^ n14490;
  assign n14495 = n14494 ^ n14486;
  assign n14496 = n14495 ^ n14488;
  assign n14497 = ~n14487 & n14496;
  assign n14498 = n14497 ^ x16;
  assign n14707 = n14706 ^ n14498;
  assign n14482 = n14460 ^ n14269;
  assign n14483 = ~n14461 & ~n14482;
  assign n14484 = n14483 ^ n14272;
  assign n14708 = n14707 ^ n14484;
  assign n14730 = n14729 ^ n14708;
  assign n14956 = n14708 & ~n14711;
  assign n14957 = ~n14480 & ~n14956;
  assign n14958 = ~n14708 & ~n14713;
  assign n14959 = ~n14712 & ~n14958;
  assign n14960 = ~n14957 & n14959;
  assign n14961 = ~n14708 & ~n14709;
  assign n14962 = n14462 ^ n14258;
  assign n14963 = n14480 ^ n14462;
  assign n14964 = ~n14962 & n14963;
  assign n14965 = n14964 ^ n14462;
  assign n14966 = ~n14961 & n14965;
  assign n14967 = ~n14960 & ~n14966;
  assign n14945 = n1404 & ~n10855;
  assign n14946 = x126 & n1408;
  assign n14947 = x125 & n1514;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = x127 & n1517;
  assign n14950 = n14948 & ~n14949;
  assign n14951 = ~n14945 & n14950;
  assign n14952 = n14951 ^ x20;
  assign n14935 = n1746 & n9999;
  assign n14936 = x123 & n1750;
  assign n14937 = x122 & n1871;
  assign n14938 = ~n14936 & ~n14937;
  assign n14939 = x124 & n1873;
  assign n14940 = n14938 & ~n14939;
  assign n14941 = ~n14935 & n14940;
  assign n14942 = n14941 ^ x23;
  assign n14923 = n2527 & n8265;
  assign n14924 = x116 & n2690;
  assign n14925 = x117 & n2530;
  assign n14926 = ~n14924 & ~n14925;
  assign n14927 = x118 & n2693;
  assign n14928 = n14926 & ~n14927;
  assign n14929 = ~n14923 & n14928;
  assign n14930 = n14929 ^ x29;
  assign n14913 = n3009 & n7481;
  assign n14914 = x113 & n3181;
  assign n14915 = x114 & n3013;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = x115 & n3183;
  assign n14918 = n14916 & ~n14917;
  assign n14919 = ~n14913 & n14918;
  assign n14920 = n14919 ^ x32;
  assign n14903 = n3522 & n6728;
  assign n14904 = x110 & n3699;
  assign n14905 = x112 & n3701;
  assign n14906 = ~n14904 & ~n14905;
  assign n14907 = x111 & n3526;
  assign n14908 = n14906 & ~n14907;
  assign n14909 = ~n14903 & n14908;
  assign n14910 = n14909 ^ x35;
  assign n14893 = n4040 & n6026;
  assign n14894 = x107 & n4267;
  assign n14895 = x108 & n4044;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = x109 & n4270;
  assign n14898 = n14896 & ~n14897;
  assign n14899 = ~n14893 & n14898;
  assign n14900 = n14899 ^ x38;
  assign n14883 = n4643 & n5351;
  assign n14884 = x104 & n4653;
  assign n14885 = x105 & n4646;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = x106 & n5046;
  assign n14888 = n14886 & ~n14887;
  assign n14889 = ~n14883 & n14888;
  assign n14890 = n14889 ^ x41;
  assign n14873 = n4718 & n5262;
  assign n14874 = x101 & n5488;
  assign n14875 = x103 & n5491;
  assign n14876 = ~n14874 & ~n14875;
  assign n14877 = x102 & n5266;
  assign n14878 = n14876 & ~n14877;
  assign n14879 = ~n14873 & n14878;
  assign n14880 = n14879 ^ x44;
  assign n14863 = n4141 & n5942;
  assign n14864 = x98 & n6186;
  assign n14865 = x99 & n5947;
  assign n14866 = ~n14864 & ~n14865;
  assign n14867 = x100 & n6406;
  assign n14868 = n14866 & ~n14867;
  assign n14869 = ~n14863 & n14868;
  assign n14870 = n14869 ^ x47;
  assign n14853 = n3585 & n6626;
  assign n14854 = x96 & n6630;
  assign n14855 = x95 & n6884;
  assign n14856 = ~n14854 & ~n14855;
  assign n14857 = x97 & n6888;
  assign n14858 = n14856 & ~n14857;
  assign n14859 = ~n14853 & n14858;
  assign n14860 = n14859 ^ x50;
  assign n14843 = n3078 & n7395;
  assign n14844 = x93 & n7400;
  assign n14845 = x92 & n7650;
  assign n14846 = ~n14844 & ~n14845;
  assign n14847 = x94 & n7652;
  assign n14848 = n14846 & ~n14847;
  assign n14849 = ~n14843 & n14848;
  assign n14850 = n14849 ^ x53;
  assign n14831 = n2176 & n9002;
  assign n14832 = x86 & n9012;
  assign n14833 = x87 & n9005;
  assign n14834 = ~n14832 & ~n14833;
  assign n14835 = x88 & n9557;
  assign n14836 = n14834 & ~n14835;
  assign n14837 = ~n14831 & n14836;
  assign n14838 = n14837 ^ x59;
  assign n14828 = n14572 ^ n14544;
  assign n14829 = n14564 & n14828;
  assign n14830 = n14829 ^ n14572;
  assign n14839 = n14838 ^ n14830;
  assign n14807 = x80 & ~x81;
  assign n14808 = x63 & n14807;
  assign n14809 = ~x62 & ~n14808;
  assign n14810 = n14562 & n14809;
  assign n14811 = n14562 ^ x81;
  assign n14812 = ~n1130 & ~n14811;
  assign n14813 = n14812 ^ x81;
  assign n14814 = n14116 & n14813;
  assign n14815 = ~n14810 & ~n14814;
  assign n14816 = ~x80 & x81;
  assign n14817 = n14816 ^ x62;
  assign n14818 = n14817 ^ n14816;
  assign n14819 = n14562 ^ x80;
  assign n14820 = ~n1030 & ~n14819;
  assign n14821 = n14820 ^ x80;
  assign n14822 = n14821 ^ n14816;
  assign n14823 = n14818 & n14822;
  assign n14824 = n14823 ^ n14816;
  assign n14825 = x63 & n14824;
  assign n14826 = n14815 & ~n14825;
  assign n14798 = n1801 & n9878;
  assign n14799 = x83 & n9888;
  assign n14800 = x85 & n10501;
  assign n14801 = ~n14799 & ~n14800;
  assign n14802 = x84 & n9881;
  assign n14803 = n14801 & ~n14802;
  assign n14804 = ~n14798 & n14803;
  assign n14805 = n14804 ^ x62;
  assign n14789 = n1225 ^ x63;
  assign n14790 = n14789 ^ n1225;
  assign n14791 = n1225 ^ n1130;
  assign n14792 = n14791 ^ n1225;
  assign n14793 = n14790 & n14792;
  assign n14794 = n14793 ^ n1225;
  assign n14795 = ~n10177 & n14794;
  assign n14796 = n14795 ^ n1225;
  assign n14797 = n14796 ^ x17;
  assign n14806 = n14805 ^ n14797;
  assign n14827 = n14826 ^ n14806;
  assign n14840 = n14839 ^ n14827;
  assign n14781 = n2607 & n8171;
  assign n14782 = x89 & n8181;
  assign n14783 = x91 & n8732;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = x90 & n8174;
  assign n14786 = n14784 & ~n14785;
  assign n14787 = ~n14781 & n14786;
  assign n14788 = n14787 ^ x56;
  assign n14841 = n14840 ^ n14788;
  assign n14778 = n14582 ^ n14534;
  assign n14779 = n14574 & n14778;
  assign n14780 = n14779 ^ n14582;
  assign n14842 = n14841 ^ n14780;
  assign n14851 = n14850 ^ n14842;
  assign n14775 = n14583 ^ n14531;
  assign n14776 = ~n14592 & n14775;
  assign n14777 = n14776 ^ n14591;
  assign n14852 = n14851 ^ n14777;
  assign n14861 = n14860 ^ n14852;
  assign n14772 = n14593 ^ n14528;
  assign n14773 = ~n14602 & n14772;
  assign n14774 = n14773 ^ n14601;
  assign n14862 = n14861 ^ n14774;
  assign n14871 = n14870 ^ n14862;
  assign n14769 = n14606 ^ n14603;
  assign n14770 = n14615 & n14769;
  assign n14771 = n14770 ^ n14614;
  assign n14872 = n14871 ^ n14771;
  assign n14881 = n14880 ^ n14872;
  assign n14766 = n14616 ^ n14525;
  assign n14767 = ~n14625 & n14766;
  assign n14768 = n14767 ^ n14624;
  assign n14882 = n14881 ^ n14768;
  assign n14891 = n14890 ^ n14882;
  assign n14763 = n14635 ^ n14522;
  assign n14764 = n14627 & n14763;
  assign n14765 = n14764 ^ n14635;
  assign n14892 = n14891 ^ n14765;
  assign n14901 = n14900 ^ n14892;
  assign n14760 = n14645 ^ n14636;
  assign n14761 = n14637 & ~n14760;
  assign n14762 = n14761 ^ n14645;
  assign n14902 = n14901 ^ n14762;
  assign n14911 = n14910 ^ n14902;
  assign n14757 = n14655 ^ n14516;
  assign n14758 = n14647 & n14757;
  assign n14759 = n14758 ^ n14655;
  assign n14912 = n14911 ^ n14759;
  assign n14921 = n14920 ^ n14912;
  assign n14754 = n14665 ^ n14656;
  assign n14755 = n14657 & ~n14754;
  assign n14756 = n14755 ^ n14665;
  assign n14922 = n14921 ^ n14756;
  assign n14931 = n14930 ^ n14922;
  assign n14751 = n14675 ^ n14666;
  assign n14752 = n14667 & ~n14751;
  assign n14753 = n14752 ^ n14675;
  assign n14932 = n14931 ^ n14753;
  assign n14748 = n14685 ^ n14676;
  assign n14749 = n14677 & ~n14748;
  assign n14750 = n14749 ^ n14685;
  assign n14933 = n14932 ^ n14750;
  assign n14740 = n2102 & n9094;
  assign n14741 = x119 & n2112;
  assign n14742 = x120 & n2105;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = x121 & n2381;
  assign n14745 = n14743 & ~n14744;
  assign n14746 = ~n14740 & n14745;
  assign n14747 = n14746 ^ x26;
  assign n14934 = n14933 ^ n14747;
  assign n14943 = n14942 ^ n14934;
  assign n14737 = n14695 ^ n14504;
  assign n14738 = ~n14687 & ~n14737;
  assign n14739 = n14738 ^ n14695;
  assign n14944 = n14943 ^ n14739;
  assign n14953 = n14952 ^ n14944;
  assign n14734 = n14705 ^ n14501;
  assign n14735 = n14697 & ~n14734;
  assign n14736 = n14735 ^ n14705;
  assign n14954 = n14953 ^ n14736;
  assign n14731 = n14498 ^ n14484;
  assign n14732 = ~n14707 & n14731;
  assign n14733 = n14732 ^ n14484;
  assign n14955 = n14954 ^ n14733;
  assign n14968 = n14967 ^ n14955;
  assign n15181 = n1746 & n10303;
  assign n15182 = x124 & n1750;
  assign n15183 = x123 & n1871;
  assign n15184 = ~n15182 & ~n15183;
  assign n15185 = x125 & n1873;
  assign n15186 = n15184 & ~n15185;
  assign n15187 = ~n15181 & n15186;
  assign n15188 = n15187 ^ x23;
  assign n15171 = n2102 & n9387;
  assign n15172 = x120 & n2112;
  assign n15173 = x121 & n2105;
  assign n15174 = ~n15172 & ~n15173;
  assign n15175 = x122 & n2381;
  assign n15176 = n15174 & ~n15175;
  assign n15177 = ~n15171 & n15176;
  assign n15178 = n15177 ^ x26;
  assign n15160 = n2527 & n8542;
  assign n15161 = x117 & n2690;
  assign n15162 = x119 & n2693;
  assign n15163 = ~n15161 & ~n15162;
  assign n15164 = x118 & n2530;
  assign n15165 = n15163 & ~n15164;
  assign n15166 = ~n15160 & n15165;
  assign n15167 = n15166 ^ x29;
  assign n15151 = n3009 & n7730;
  assign n15152 = x114 & n3181;
  assign n15153 = x115 & n3013;
  assign n15154 = ~n15152 & ~n15153;
  assign n15155 = x116 & n3183;
  assign n15156 = n15154 & ~n15155;
  assign n15157 = ~n15151 & n15156;
  assign n15158 = n15157 ^ x32;
  assign n15141 = n3522 & n6975;
  assign n15142 = x111 & n3699;
  assign n15143 = x113 & n3701;
  assign n15144 = ~n15142 & ~n15143;
  assign n15145 = x112 & n3526;
  assign n15146 = n15144 & ~n15145;
  assign n15147 = ~n15141 & n15146;
  assign n15148 = n15147 ^ x35;
  assign n15125 = n4323 & n5942;
  assign n15126 = x99 & n6186;
  assign n15127 = x101 & n6406;
  assign n15128 = ~n15126 & ~n15127;
  assign n15129 = x100 & n5947;
  assign n15130 = n15128 & ~n15129;
  assign n15131 = ~n15125 & n15130;
  assign n15132 = n15131 ^ x47;
  assign n15115 = n3763 & n6626;
  assign n15116 = x96 & n6884;
  assign n15117 = x98 & n6888;
  assign n15118 = ~n15116 & ~n15117;
  assign n15119 = x97 & n6630;
  assign n15120 = n15118 & ~n15119;
  assign n15121 = ~n15115 & n15120;
  assign n15122 = n15121 ^ x50;
  assign n15105 = n3247 & n7395;
  assign n15106 = x93 & n7650;
  assign n15107 = x94 & n7400;
  assign n15108 = ~n15106 & ~n15107;
  assign n15109 = x95 & n7652;
  assign n15110 = n15108 & ~n15109;
  assign n15111 = ~n15105 & n15110;
  assign n15112 = n15111 ^ x53;
  assign n15094 = n2755 & n8171;
  assign n15095 = x90 & n8181;
  assign n15096 = x91 & n8174;
  assign n15097 = ~n15095 & ~n15096;
  assign n15098 = x92 & n8732;
  assign n15099 = n15097 & ~n15098;
  assign n15100 = ~n15094 & n15099;
  assign n15101 = n15100 ^ x56;
  assign n15091 = n14838 ^ n14827;
  assign n15092 = n14839 & n15091;
  assign n15093 = n15092 ^ n14830;
  assign n15102 = n15101 ^ n15093;
  assign n15081 = n2310 & n9002;
  assign n15082 = x88 & n9005;
  assign n15083 = x89 & n9557;
  assign n15084 = ~n15082 & ~n15083;
  assign n15085 = x87 & n9012;
  assign n15086 = n15084 & ~n15085;
  assign n15087 = ~n15081 & n15086;
  assign n15088 = n15087 ^ x59;
  assign n15072 = n1920 & n9878;
  assign n15073 = x84 & n9888;
  assign n15074 = x85 & n9881;
  assign n15075 = ~n15073 & ~n15074;
  assign n15076 = x86 & n10501;
  assign n15077 = n15075 & ~n15076;
  assign n15078 = ~n15072 & n15077;
  assign n15079 = n15078 ^ x62;
  assign n15068 = x83 & n10177;
  assign n15069 = x82 & n12123;
  assign n15070 = ~n15068 & ~n15069;
  assign n15058 = x81 ^ x17;
  assign n15059 = x82 ^ x80;
  assign n15060 = n12123 ^ x82;
  assign n15061 = n15060 ^ x82;
  assign n15062 = n15059 & n15061;
  assign n15063 = n15062 ^ x82;
  assign n15064 = n15063 ^ x81;
  assign n15065 = ~n15058 & n15064;
  assign n15066 = n15065 ^ x81;
  assign n15067 = ~n12893 & n15066;
  assign n15071 = n15070 ^ n15067;
  assign n15080 = n15079 ^ n15071;
  assign n15089 = n15088 ^ n15080;
  assign n15055 = n14826 ^ n14805;
  assign n15056 = ~n14806 & ~n15055;
  assign n15057 = n15056 ^ n14826;
  assign n15090 = n15089 ^ n15057;
  assign n15103 = n15102 ^ n15090;
  assign n15052 = n14788 ^ n14780;
  assign n15053 = ~n14841 & ~n15052;
  assign n15054 = n15053 ^ n14840;
  assign n15104 = n15103 ^ n15054;
  assign n15113 = n15112 ^ n15104;
  assign n15049 = n14850 ^ n14777;
  assign n15050 = n14851 & n15049;
  assign n15051 = n15050 ^ n14777;
  assign n15114 = n15113 ^ n15051;
  assign n15123 = n15122 ^ n15114;
  assign n15046 = n14860 ^ n14774;
  assign n15047 = n14861 & n15046;
  assign n15048 = n15047 ^ n14774;
  assign n15124 = n15123 ^ n15048;
  assign n15133 = n15132 ^ n15124;
  assign n15043 = n14870 ^ n14771;
  assign n15044 = n14871 & n15043;
  assign n15045 = n15044 ^ n14771;
  assign n15134 = n15133 ^ n15045;
  assign n15035 = n4912 & n5262;
  assign n15036 = x102 & n5488;
  assign n15037 = x103 & n5266;
  assign n15038 = ~n15036 & ~n15037;
  assign n15039 = x104 & n5491;
  assign n15040 = n15038 & ~n15039;
  assign n15041 = ~n15035 & n15040;
  assign n15042 = n15041 ^ x44;
  assign n15135 = n15134 ^ n15042;
  assign n15032 = n14880 ^ n14768;
  assign n15033 = n14881 & n15032;
  assign n15034 = n15033 ^ n14768;
  assign n15136 = n15135 ^ n15034;
  assign n15024 = n4643 & n5578;
  assign n15025 = x105 & n4653;
  assign n15026 = x107 & n5046;
  assign n15027 = ~n15025 & ~n15026;
  assign n15028 = x106 & n4646;
  assign n15029 = n15027 & ~n15028;
  assign n15030 = ~n15024 & n15029;
  assign n15031 = n15030 ^ x41;
  assign n15137 = n15136 ^ n15031;
  assign n15021 = n14890 ^ n14765;
  assign n15022 = n14891 & n15021;
  assign n15023 = n15022 ^ n14765;
  assign n15138 = n15137 ^ n15023;
  assign n15013 = n4040 & n6250;
  assign n15014 = x108 & n4267;
  assign n15015 = x109 & n4044;
  assign n15016 = ~n15014 & ~n15015;
  assign n15017 = x110 & n4270;
  assign n15018 = n15016 & ~n15017;
  assign n15019 = ~n15013 & n15018;
  assign n15020 = n15019 ^ x38;
  assign n15139 = n15138 ^ n15020;
  assign n15010 = n14900 ^ n14762;
  assign n15011 = n14901 & n15010;
  assign n15012 = n15011 ^ n14762;
  assign n15140 = n15139 ^ n15012;
  assign n15149 = n15148 ^ n15140;
  assign n15007 = n14902 ^ n14759;
  assign n15008 = ~n14911 & n15007;
  assign n15009 = n15008 ^ n14910;
  assign n15150 = n15149 ^ n15009;
  assign n15159 = n15158 ^ n15150;
  assign n15168 = n15167 ^ n15159;
  assign n15004 = n14920 ^ n14756;
  assign n15005 = n14921 & n15004;
  assign n15006 = n15005 ^ n14756;
  assign n15169 = n15168 ^ n15006;
  assign n15001 = n14930 ^ n14753;
  assign n15002 = n14931 & n15001;
  assign n15003 = n15002 ^ n14753;
  assign n15170 = n15169 ^ n15003;
  assign n15179 = n15178 ^ n15170;
  assign n14998 = n14932 ^ n14747;
  assign n14999 = ~n14933 & n14998;
  assign n15000 = n14999 ^ n14750;
  assign n15180 = n15179 ^ n15000;
  assign n15189 = n15188 ^ n15180;
  assign n14995 = n14942 ^ n14739;
  assign n14996 = n14943 & n14995;
  assign n14997 = n14996 ^ n14739;
  assign n15190 = n15189 ^ n14997;
  assign n14989 = n1404 & ~n10281;
  assign n14990 = x127 & n1408;
  assign n14991 = x126 & n1514;
  assign n14992 = ~n14990 & ~n14991;
  assign n14993 = ~n14989 & n14992;
  assign n14994 = n14993 ^ x20;
  assign n15191 = n15190 ^ n14994;
  assign n14969 = n14733 & ~n14736;
  assign n14970 = ~n14952 & n14969;
  assign n14971 = ~n14733 & n14736;
  assign n14972 = n14952 & n14971;
  assign n14973 = ~n14970 & ~n14972;
  assign n14974 = n14953 & ~n14973;
  assign n14975 = ~n14944 & ~n14970;
  assign n14976 = n14952 ^ n14733;
  assign n14977 = n14952 ^ n14736;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = n14978 ^ n14733;
  assign n14980 = ~n14975 & n14979;
  assign n14981 = n14980 ^ n14967;
  assign n14982 = n14981 ^ n14980;
  assign n14983 = n14944 & ~n14972;
  assign n14984 = ~n14979 & ~n14983;
  assign n14985 = n14984 ^ n14980;
  assign n14986 = n14982 & n14985;
  assign n14987 = n14986 ^ n14980;
  assign n14988 = ~n14974 & ~n14987;
  assign n15192 = n15191 ^ n14988;
  assign n15414 = n14944 & ~n14952;
  assign n15415 = ~n14971 & n15414;
  assign n15416 = n15191 & ~n15415;
  assign n15417 = ~n14967 & ~n15416;
  assign n15418 = ~n14944 & n14952;
  assign n15419 = ~n15191 & ~n15418;
  assign n15420 = ~n14969 & ~n15419;
  assign n15421 = ~n15417 & n15420;
  assign n15422 = ~n14971 & ~n15191;
  assign n15423 = n14967 ^ n14952;
  assign n15424 = ~n14953 & n15423;
  assign n15425 = n15424 ^ n14952;
  assign n15426 = ~n15422 & n15425;
  assign n15427 = ~n15421 & ~n15426;
  assign n15403 = n1746 & ~n10570;
  assign n15404 = x124 & n1871;
  assign n15405 = x125 & n1750;
  assign n15406 = ~n15404 & ~n15405;
  assign n15407 = x126 & n1873;
  assign n15408 = n15406 & ~n15407;
  assign n15409 = ~n15403 & n15408;
  assign n15410 = n15409 ^ x23;
  assign n15393 = n2102 & n9691;
  assign n15394 = x121 & n2112;
  assign n15395 = x122 & n2105;
  assign n15396 = ~n15394 & ~n15395;
  assign n15397 = x123 & n2381;
  assign n15398 = n15396 & ~n15397;
  assign n15399 = ~n15393 & n15398;
  assign n15400 = n15399 ^ x26;
  assign n15383 = n2527 & n8820;
  assign n15384 = x118 & n2690;
  assign n15385 = x119 & n2530;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = x120 & n2693;
  assign n15388 = n15386 & ~n15387;
  assign n15389 = ~n15383 & n15388;
  assign n15390 = n15389 ^ x29;
  assign n15373 = n3009 & n7987;
  assign n15374 = x116 & n3013;
  assign n15375 = x115 & n3181;
  assign n15376 = ~n15374 & ~n15375;
  assign n15377 = x117 & n3183;
  assign n15378 = n15376 & ~n15377;
  assign n15379 = ~n15373 & n15378;
  assign n15380 = n15379 ^ x32;
  assign n15363 = n3522 & n7220;
  assign n15364 = x112 & n3699;
  assign n15365 = x114 & n3701;
  assign n15366 = ~n15364 & ~n15365;
  assign n15367 = x113 & n3526;
  assign n15368 = n15366 & ~n15367;
  assign n15369 = ~n15363 & n15368;
  assign n15370 = n15369 ^ x35;
  assign n15353 = n4040 & n6478;
  assign n15354 = x109 & n4267;
  assign n15355 = x111 & n4270;
  assign n15356 = ~n15354 & ~n15355;
  assign n15357 = x110 & n4044;
  assign n15358 = n15356 & ~n15357;
  assign n15359 = ~n15353 & n15358;
  assign n15360 = n15359 ^ x38;
  assign n15343 = n4643 & n5792;
  assign n15344 = x106 & n4653;
  assign n15345 = x108 & n5046;
  assign n15346 = ~n15344 & ~n15345;
  assign n15347 = x107 & n4646;
  assign n15348 = n15346 & ~n15347;
  assign n15349 = ~n15343 & n15348;
  assign n15350 = n15349 ^ x41;
  assign n15333 = n5117 & n5262;
  assign n15334 = x103 & n5488;
  assign n15335 = x104 & n5266;
  assign n15336 = ~n15334 & ~n15335;
  assign n15337 = x105 & n5491;
  assign n15338 = n15336 & ~n15337;
  assign n15339 = ~n15333 & n15338;
  assign n15340 = n15339 ^ x44;
  assign n15320 = n3943 & n6626;
  assign n15321 = x97 & n6884;
  assign n15322 = x99 & n6888;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = x98 & n6630;
  assign n15325 = n15323 & ~n15324;
  assign n15326 = ~n15320 & n15325;
  assign n15327 = n15326 ^ x50;
  assign n15317 = n15112 ^ n15054;
  assign n15318 = ~n15104 & ~n15317;
  assign n15319 = n15318 ^ n15112;
  assign n15328 = n15327 ^ n15319;
  assign n15307 = n3403 & n7395;
  assign n15308 = x94 & n7650;
  assign n15309 = x96 & n7652;
  assign n15310 = ~n15308 & ~n15309;
  assign n15311 = x95 & n7400;
  assign n15312 = n15310 & ~n15311;
  assign n15313 = ~n15307 & n15312;
  assign n15314 = n15313 ^ x53;
  assign n15297 = n2901 & n8171;
  assign n15298 = x91 & n8181;
  assign n15299 = x92 & n8174;
  assign n15300 = ~n15298 & ~n15299;
  assign n15301 = x93 & n8732;
  assign n15302 = n15300 & ~n15301;
  assign n15303 = ~n15297 & n15302;
  assign n15304 = n15303 ^ x56;
  assign n15294 = n15080 ^ n15057;
  assign n15295 = n15089 & n15294;
  assign n15296 = n15295 ^ n15088;
  assign n15305 = n15304 ^ n15296;
  assign n15285 = n2448 & n9002;
  assign n15286 = x88 & n9012;
  assign n15287 = x89 & n9005;
  assign n15288 = ~n15286 & ~n15287;
  assign n15289 = x90 & n9557;
  assign n15290 = n15288 & ~n15289;
  assign n15291 = ~n15285 & n15290;
  assign n15292 = n15291 ^ x59;
  assign n15275 = n2039 & n9878;
  assign n15276 = x85 & n9888;
  assign n15277 = x86 & n9881;
  assign n15278 = ~n15276 & ~n15277;
  assign n15279 = x87 & n10501;
  assign n15280 = n15278 & ~n15279;
  assign n15281 = ~n15275 & n15280;
  assign n15282 = n15281 ^ x62;
  assign n15255 = n15069 ^ x84;
  assign n15256 = n15255 ^ n15069;
  assign n15257 = n15069 ^ n10177;
  assign n15258 = n15257 ^ n15069;
  assign n15259 = ~n15256 & n15258;
  assign n15260 = n15259 ^ n15069;
  assign n15261 = x83 & n15260;
  assign n15262 = n15261 ^ n15069;
  assign n15263 = n10177 ^ x83;
  assign n15264 = n1443 ^ x84;
  assign n15265 = n15264 ^ n15263;
  assign n15266 = x82 ^ x63;
  assign n15267 = ~x82 & ~n15266;
  assign n15268 = n15267 ^ x84;
  assign n15269 = n15268 ^ x82;
  assign n15270 = n15265 & ~n15269;
  assign n15271 = n15270 ^ n15267;
  assign n15272 = n15271 ^ x82;
  assign n15273 = n15263 & ~n15272;
  assign n15274 = ~n15262 & ~n15273;
  assign n15283 = n15282 ^ n15274;
  assign n15252 = n15079 ^ n15067;
  assign n15253 = ~n15071 & ~n15252;
  assign n15254 = n15253 ^ n15079;
  assign n15284 = n15283 ^ n15254;
  assign n15293 = n15292 ^ n15284;
  assign n15306 = n15305 ^ n15293;
  assign n15315 = n15314 ^ n15306;
  assign n15249 = n15101 ^ n15090;
  assign n15250 = n15102 & n15249;
  assign n15251 = n15250 ^ n15093;
  assign n15316 = n15315 ^ n15251;
  assign n15329 = n15328 ^ n15316;
  assign n15246 = n15122 ^ n15051;
  assign n15247 = ~n15114 & n15246;
  assign n15248 = n15247 ^ n15122;
  assign n15330 = n15329 ^ n15248;
  assign n15238 = n4509 & n5942;
  assign n15239 = x101 & n5947;
  assign n15240 = x100 & n6186;
  assign n15241 = ~n15239 & ~n15240;
  assign n15242 = x102 & n6406;
  assign n15243 = n15241 & ~n15242;
  assign n15244 = ~n15238 & n15243;
  assign n15245 = n15244 ^ x47;
  assign n15331 = n15330 ^ n15245;
  assign n15235 = n15132 ^ n15048;
  assign n15236 = ~n15124 & n15235;
  assign n15237 = n15236 ^ n15132;
  assign n15332 = n15331 ^ n15237;
  assign n15341 = n15340 ^ n15332;
  assign n15232 = n15133 ^ n15042;
  assign n15233 = n15134 & ~n15232;
  assign n15234 = n15233 ^ n15045;
  assign n15342 = n15341 ^ n15234;
  assign n15351 = n15350 ^ n15342;
  assign n15229 = n15135 ^ n15031;
  assign n15230 = n15136 & ~n15229;
  assign n15231 = n15230 ^ n15034;
  assign n15352 = n15351 ^ n15231;
  assign n15361 = n15360 ^ n15352;
  assign n15226 = n15137 ^ n15020;
  assign n15227 = n15138 & ~n15226;
  assign n15228 = n15227 ^ n15023;
  assign n15362 = n15361 ^ n15228;
  assign n15371 = n15370 ^ n15362;
  assign n15223 = n15148 ^ n15139;
  assign n15224 = ~n15140 & n15223;
  assign n15225 = n15224 ^ n15148;
  assign n15372 = n15371 ^ n15225;
  assign n15381 = n15380 ^ n15372;
  assign n15220 = n15158 ^ n15009;
  assign n15221 = ~n15150 & n15220;
  assign n15222 = n15221 ^ n15158;
  assign n15382 = n15381 ^ n15222;
  assign n15391 = n15390 ^ n15382;
  assign n15217 = n15159 ^ n15006;
  assign n15218 = n15168 & ~n15217;
  assign n15219 = n15218 ^ n15167;
  assign n15392 = n15391 ^ n15219;
  assign n15401 = n15400 ^ n15392;
  assign n15214 = n15178 ^ n15003;
  assign n15215 = ~n15170 & n15214;
  assign n15216 = n15215 ^ n15178;
  assign n15402 = n15401 ^ n15216;
  assign n15411 = n15410 ^ n15402;
  assign n15211 = n15189 ^ n14994;
  assign n15212 = n15190 & ~n15211;
  assign n15213 = n15212 ^ n14997;
  assign n15412 = n15411 ^ n15213;
  assign n15196 = x127 & n1284;
  assign n15197 = ~x20 & ~n15196;
  assign n15198 = n15197 ^ x19;
  assign n15199 = n1191 & n11409;
  assign n15200 = n15199 ^ n15197;
  assign n15201 = ~n15197 & n15200;
  assign n15202 = n15201 ^ n15197;
  assign n15203 = x127 & n1513;
  assign n15204 = ~n15202 & ~n15203;
  assign n15205 = n15204 ^ n15201;
  assign n15206 = n15205 ^ n15197;
  assign n15207 = n15206 ^ n15199;
  assign n15208 = ~n15198 & n15207;
  assign n15209 = n15208 ^ x19;
  assign n15193 = n15188 ^ n15179;
  assign n15194 = ~n15180 & n15193;
  assign n15195 = n15194 ^ n15188;
  assign n15210 = n15209 ^ n15195;
  assign n15413 = n15412 ^ n15210;
  assign n15428 = n15427 ^ n15413;
  assign n15620 = ~n15195 & n15209;
  assign n15625 = n15213 & n15411;
  assign n15626 = ~n15620 & n15625;
  assign n15619 = n15195 & ~n15209;
  assign n15627 = ~n15213 & ~n15411;
  assign n15628 = n15619 & ~n15627;
  assign n15629 = ~n15626 & ~n15628;
  assign n15621 = n15620 ^ n15411;
  assign n15622 = n15412 & n15621;
  assign n15623 = n15622 ^ n15213;
  assign n15624 = ~n15619 & ~n15623;
  assign n15630 = n15629 ^ n15624;
  assign n15631 = n15427 & ~n15630;
  assign n15632 = n15631 ^ n15629;
  assign n15633 = n15411 ^ n15209;
  assign n15634 = n15210 & n15633;
  assign n15635 = ~n15412 & n15634;
  assign n15636 = n15632 & ~n15635;
  assign n15609 = n1746 & ~n10855;
  assign n15610 = x126 & n1750;
  assign n15611 = x125 & n1871;
  assign n15612 = ~n15610 & ~n15611;
  assign n15613 = x127 & n1873;
  assign n15614 = n15612 & ~n15613;
  assign n15615 = ~n15609 & n15614;
  assign n15616 = n15615 ^ x23;
  assign n15599 = n2102 & n9999;
  assign n15600 = x122 & n2112;
  assign n15601 = x123 & n2105;
  assign n15602 = ~n15600 & ~n15601;
  assign n15603 = x124 & n2381;
  assign n15604 = n15602 & ~n15603;
  assign n15605 = ~n15599 & n15604;
  assign n15606 = n15605 ^ x26;
  assign n15587 = n3009 & n8265;
  assign n15588 = x116 & n3181;
  assign n15589 = x117 & n3013;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = x118 & n3183;
  assign n15592 = n15590 & ~n15591;
  assign n15593 = ~n15587 & n15592;
  assign n15594 = n15593 ^ x32;
  assign n15577 = n3522 & n7481;
  assign n15578 = x113 & n3699;
  assign n15579 = x114 & n3526;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = x115 & n3701;
  assign n15582 = n15580 & ~n15581;
  assign n15583 = ~n15577 & n15582;
  assign n15584 = n15583 ^ x35;
  assign n15567 = n4040 & n6728;
  assign n15568 = x110 & n4267;
  assign n15569 = x112 & n4270;
  assign n15570 = ~n15568 & ~n15569;
  assign n15571 = x111 & n4044;
  assign n15572 = n15570 & ~n15571;
  assign n15573 = ~n15567 & n15572;
  assign n15574 = n15573 ^ x38;
  assign n15557 = n4643 & n6026;
  assign n15558 = x107 & n4653;
  assign n15559 = x108 & n4646;
  assign n15560 = ~n15558 & ~n15559;
  assign n15561 = x109 & n5046;
  assign n15562 = n15560 & ~n15561;
  assign n15563 = ~n15557 & n15562;
  assign n15564 = n15563 ^ x41;
  assign n15547 = n5262 & n5351;
  assign n15548 = x105 & n5266;
  assign n15549 = x104 & n5488;
  assign n15550 = ~n15548 & ~n15549;
  assign n15551 = x106 & n5491;
  assign n15552 = n15550 & ~n15551;
  assign n15553 = ~n15547 & n15552;
  assign n15554 = n15553 ^ x44;
  assign n15535 = n4141 & n6626;
  assign n15536 = x98 & n6884;
  assign n15537 = x100 & n6888;
  assign n15538 = ~n15536 & ~n15537;
  assign n15539 = x99 & n6630;
  assign n15540 = n15538 & ~n15539;
  assign n15541 = ~n15535 & n15540;
  assign n15542 = n15541 ^ x50;
  assign n15532 = n15319 ^ n15316;
  assign n15533 = n15328 & ~n15532;
  assign n15534 = n15533 ^ n15327;
  assign n15543 = n15542 ^ n15534;
  assign n15522 = n3585 & n7395;
  assign n15523 = x95 & n7650;
  assign n15524 = x96 & n7400;
  assign n15525 = ~n15523 & ~n15524;
  assign n15526 = x97 & n7652;
  assign n15527 = n15525 & ~n15526;
  assign n15528 = ~n15522 & n15527;
  assign n15529 = n15528 ^ x53;
  assign n15512 = n3078 & n8171;
  assign n15513 = x92 & n8181;
  assign n15514 = x93 & n8174;
  assign n15515 = ~n15513 & ~n15514;
  assign n15516 = x94 & n8732;
  assign n15517 = n15515 & ~n15516;
  assign n15518 = ~n15512 & n15517;
  assign n15519 = n15518 ^ x56;
  assign n15502 = n2607 & n9002;
  assign n15503 = x89 & n9012;
  assign n15504 = x90 & n9005;
  assign n15505 = ~n15503 & ~n15504;
  assign n15506 = x91 & n9557;
  assign n15507 = n15505 & ~n15506;
  assign n15508 = ~n15502 & n15507;
  assign n15509 = n15508 ^ x59;
  assign n15499 = n15292 ^ n15254;
  assign n15500 = ~n15284 & n15499;
  assign n15501 = n15500 ^ n15292;
  assign n15510 = n15509 ^ n15501;
  assign n15489 = n2176 & n9878;
  assign n15490 = x86 & n9888;
  assign n15491 = x88 & n10501;
  assign n15492 = ~n15490 & ~n15491;
  assign n15493 = x87 & n9881;
  assign n15494 = n15492 & ~n15493;
  assign n15495 = ~n15489 & n15494;
  assign n15496 = n15495 ^ x62;
  assign n15480 = n1549 ^ x63;
  assign n15481 = n15480 ^ n1549;
  assign n15482 = n1549 ^ n1443;
  assign n15483 = n15482 ^ n1549;
  assign n15484 = n15481 & n15483;
  assign n15485 = n15484 ^ n1549;
  assign n15486 = ~n10177 & n15485;
  assign n15487 = n15486 ^ n1549;
  assign n15488 = n15487 ^ x20;
  assign n15497 = n15496 ^ n15488;
  assign n15478 = n15274 & ~n15282;
  assign n15479 = n15478 ^ n15262;
  assign n15498 = n15497 ^ n15479;
  assign n15511 = n15510 ^ n15498;
  assign n15520 = n15519 ^ n15511;
  assign n15475 = n15296 ^ n15293;
  assign n15476 = n15305 & ~n15475;
  assign n15477 = n15476 ^ n15304;
  assign n15521 = n15520 ^ n15477;
  assign n15530 = n15529 ^ n15521;
  assign n15472 = n15306 ^ n15251;
  assign n15473 = n15315 & ~n15472;
  assign n15474 = n15473 ^ n15314;
  assign n15531 = n15530 ^ n15474;
  assign n15544 = n15543 ^ n15531;
  assign n15469 = n15248 ^ n15245;
  assign n15470 = n15330 & ~n15469;
  assign n15471 = n15470 ^ n15329;
  assign n15545 = n15544 ^ n15471;
  assign n15461 = n4718 & n5942;
  assign n15462 = x101 & n6186;
  assign n15463 = x103 & n6406;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = x102 & n5947;
  assign n15466 = n15464 & ~n15465;
  assign n15467 = ~n15461 & n15466;
  assign n15468 = n15467 ^ x47;
  assign n15546 = n15545 ^ n15468;
  assign n15555 = n15554 ^ n15546;
  assign n15458 = n15340 ^ n15331;
  assign n15459 = ~n15332 & n15458;
  assign n15460 = n15459 ^ n15340;
  assign n15556 = n15555 ^ n15460;
  assign n15565 = n15564 ^ n15556;
  assign n15455 = n15350 ^ n15234;
  assign n15456 = ~n15342 & n15455;
  assign n15457 = n15456 ^ n15350;
  assign n15566 = n15565 ^ n15457;
  assign n15575 = n15574 ^ n15566;
  assign n15452 = n15360 ^ n15231;
  assign n15453 = ~n15352 & n15452;
  assign n15454 = n15453 ^ n15360;
  assign n15576 = n15575 ^ n15454;
  assign n15585 = n15584 ^ n15576;
  assign n15449 = n15370 ^ n15361;
  assign n15450 = ~n15362 & n15449;
  assign n15451 = n15450 ^ n15370;
  assign n15586 = n15585 ^ n15451;
  assign n15595 = n15594 ^ n15586;
  assign n15446 = n15380 ^ n15371;
  assign n15447 = ~n15372 & n15446;
  assign n15448 = n15447 ^ n15380;
  assign n15596 = n15595 ^ n15448;
  assign n15443 = n15390 ^ n15381;
  assign n15444 = ~n15382 & n15443;
  assign n15445 = n15444 ^ n15390;
  assign n15597 = n15596 ^ n15445;
  assign n15435 = n2527 & n9094;
  assign n15436 = x120 & n2530;
  assign n15437 = x119 & n2690;
  assign n15438 = ~n15436 & ~n15437;
  assign n15439 = x121 & n2693;
  assign n15440 = n15438 & ~n15439;
  assign n15441 = ~n15435 & n15440;
  assign n15442 = n15441 ^ x29;
  assign n15598 = n15597 ^ n15442;
  assign n15607 = n15606 ^ n15598;
  assign n15432 = n15400 ^ n15219;
  assign n15433 = ~n15392 & n15432;
  assign n15434 = n15433 ^ n15400;
  assign n15608 = n15607 ^ n15434;
  assign n15617 = n15616 ^ n15608;
  assign n15429 = n15410 ^ n15401;
  assign n15430 = ~n15402 & n15429;
  assign n15431 = n15430 ^ n15410;
  assign n15618 = n15617 ^ n15431;
  assign n15637 = n15636 ^ n15618;
  assign n15832 = n15618 & ~n15625;
  assign n15833 = ~n15620 & ~n15832;
  assign n15834 = n15618 & ~n15619;
  assign n15835 = ~n15627 & ~n15834;
  assign n15836 = ~n15833 & ~n15835;
  assign n15837 = ~n15427 & ~n15836;
  assign n15838 = ~n15618 & n15623;
  assign n15839 = n15619 & n15833;
  assign n15840 = ~n15838 & ~n15839;
  assign n15841 = ~n15837 & n15840;
  assign n15820 = n2102 & n10303;
  assign n15821 = x123 & n2112;
  assign n15822 = x125 & n2381;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = x124 & n2105;
  assign n15825 = n15823 & ~n15824;
  assign n15826 = ~n15820 & n15825;
  assign n15827 = n15826 ^ x26;
  assign n15810 = n2527 & n9387;
  assign n15811 = x120 & n2690;
  assign n15812 = x121 & n2530;
  assign n15813 = ~n15811 & ~n15812;
  assign n15814 = x122 & n2693;
  assign n15815 = n15813 & ~n15814;
  assign n15816 = ~n15810 & n15815;
  assign n15817 = n15816 ^ x29;
  assign n15798 = n3522 & n7730;
  assign n15799 = x114 & n3699;
  assign n15800 = x116 & n3701;
  assign n15801 = ~n15799 & ~n15800;
  assign n15802 = x115 & n3526;
  assign n15803 = n15801 & ~n15802;
  assign n15804 = ~n15798 & n15803;
  assign n15805 = n15804 ^ x35;
  assign n15788 = n4040 & n6975;
  assign n15789 = x111 & n4267;
  assign n15790 = x113 & n4270;
  assign n15791 = ~n15789 & ~n15790;
  assign n15792 = x112 & n4044;
  assign n15793 = n15791 & ~n15792;
  assign n15794 = ~n15788 & n15793;
  assign n15795 = n15794 ^ x38;
  assign n15777 = n4643 & n6250;
  assign n15778 = x108 & n4653;
  assign n15779 = x110 & n5046;
  assign n15780 = ~n15778 & ~n15779;
  assign n15781 = x109 & n4646;
  assign n15782 = n15780 & ~n15781;
  assign n15783 = ~n15777 & n15782;
  assign n15784 = n15783 ^ x41;
  assign n15768 = n5262 & n5578;
  assign n15769 = x105 & n5488;
  assign n15770 = x106 & n5266;
  assign n15771 = ~n15769 & ~n15770;
  assign n15772 = x107 & n5491;
  assign n15773 = n15771 & ~n15772;
  assign n15774 = ~n15768 & n15773;
  assign n15775 = n15774 ^ x44;
  assign n15757 = n4912 & n5942;
  assign n15758 = x102 & n6186;
  assign n15759 = x103 & n5947;
  assign n15760 = ~n15758 & ~n15759;
  assign n15761 = x104 & n6406;
  assign n15762 = n15760 & ~n15761;
  assign n15763 = ~n15757 & n15762;
  assign n15764 = n15763 ^ x47;
  assign n15754 = n15542 ^ n15531;
  assign n15755 = n15543 & n15754;
  assign n15756 = n15755 ^ n15534;
  assign n15765 = n15764 ^ n15756;
  assign n15744 = n4323 & n6626;
  assign n15745 = x99 & n6884;
  assign n15746 = x100 & n6630;
  assign n15747 = ~n15745 & ~n15746;
  assign n15748 = x101 & n6888;
  assign n15749 = n15747 & ~n15748;
  assign n15750 = ~n15744 & n15749;
  assign n15751 = n15750 ^ x50;
  assign n15734 = n3763 & n7395;
  assign n15735 = x96 & n7650;
  assign n15736 = x97 & n7400;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = x98 & n7652;
  assign n15739 = n15737 & ~n15738;
  assign n15740 = ~n15734 & n15739;
  assign n15741 = n15740 ^ x53;
  assign n15724 = n3247 & n8171;
  assign n15725 = x93 & n8181;
  assign n15726 = x95 & n8732;
  assign n15727 = ~n15725 & ~n15726;
  assign n15728 = x94 & n8174;
  assign n15729 = n15727 & ~n15728;
  assign n15730 = ~n15724 & n15729;
  assign n15731 = n15730 ^ x56;
  assign n15714 = n2755 & n9002;
  assign n15715 = x90 & n9012;
  assign n15716 = x91 & n9005;
  assign n15717 = ~n15715 & ~n15716;
  assign n15718 = x92 & n9557;
  assign n15719 = n15717 & ~n15718;
  assign n15720 = ~n15714 & n15719;
  assign n15721 = n15720 ^ x59;
  assign n15704 = n2310 & n9878;
  assign n15705 = x87 & n9888;
  assign n15706 = x89 & n10501;
  assign n15707 = ~n15705 & ~n15706;
  assign n15708 = x88 & n9881;
  assign n15709 = n15707 & ~n15708;
  assign n15710 = ~n15704 & n15709;
  assign n15711 = n15710 ^ x62;
  assign n15694 = x84 ^ x20;
  assign n15695 = x85 ^ x83;
  assign n15696 = n12123 ^ x85;
  assign n15697 = n15696 ^ x85;
  assign n15698 = n15695 & n15697;
  assign n15699 = n15698 ^ x85;
  assign n15700 = n15699 ^ x84;
  assign n15701 = ~n15694 & n15700;
  assign n15702 = n15701 ^ x84;
  assign n15703 = ~n12893 & n15702;
  assign n15712 = n15711 ^ n15703;
  assign n15691 = x86 & n10177;
  assign n15692 = x85 & n12123;
  assign n15693 = ~n15691 & ~n15692;
  assign n15713 = n15712 ^ n15693;
  assign n15722 = n15721 ^ n15713;
  assign n15688 = n15496 ^ n15479;
  assign n15689 = ~n15497 & ~n15688;
  assign n15690 = n15689 ^ n15479;
  assign n15723 = n15722 ^ n15690;
  assign n15732 = n15731 ^ n15723;
  assign n15685 = n15509 ^ n15498;
  assign n15686 = n15510 & n15685;
  assign n15687 = n15686 ^ n15501;
  assign n15733 = n15732 ^ n15687;
  assign n15742 = n15741 ^ n15733;
  assign n15682 = n15519 ^ n15477;
  assign n15683 = n15520 & n15682;
  assign n15684 = n15683 ^ n15477;
  assign n15743 = n15742 ^ n15684;
  assign n15752 = n15751 ^ n15743;
  assign n15679 = n15529 ^ n15474;
  assign n15680 = n15530 & n15679;
  assign n15681 = n15680 ^ n15474;
  assign n15753 = n15752 ^ n15681;
  assign n15766 = n15765 ^ n15753;
  assign n15676 = n15544 ^ n15468;
  assign n15677 = ~n15545 & n15676;
  assign n15678 = n15677 ^ n15471;
  assign n15767 = n15766 ^ n15678;
  assign n15776 = n15775 ^ n15767;
  assign n15785 = n15784 ^ n15776;
  assign n15673 = n15554 ^ n15460;
  assign n15674 = n15555 & n15673;
  assign n15675 = n15674 ^ n15460;
  assign n15786 = n15785 ^ n15675;
  assign n15670 = n15556 ^ n15457;
  assign n15671 = ~n15565 & n15670;
  assign n15672 = n15671 ^ n15564;
  assign n15787 = n15786 ^ n15672;
  assign n15796 = n15795 ^ n15787;
  assign n15667 = n15566 ^ n15454;
  assign n15668 = ~n15575 & n15667;
  assign n15669 = n15668 ^ n15574;
  assign n15797 = n15796 ^ n15669;
  assign n15806 = n15805 ^ n15797;
  assign n15664 = n15584 ^ n15451;
  assign n15665 = n15585 & n15664;
  assign n15666 = n15665 ^ n15451;
  assign n15807 = n15806 ^ n15666;
  assign n15656 = n3009 & n8542;
  assign n15657 = x117 & n3181;
  assign n15658 = x118 & n3013;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = x119 & n3183;
  assign n15661 = n15659 & ~n15660;
  assign n15662 = ~n15656 & n15661;
  assign n15663 = n15662 ^ x32;
  assign n15808 = n15807 ^ n15663;
  assign n15653 = n15594 ^ n15448;
  assign n15654 = n15595 & n15653;
  assign n15655 = n15654 ^ n15448;
  assign n15809 = n15808 ^ n15655;
  assign n15818 = n15817 ^ n15809;
  assign n15650 = n15596 ^ n15442;
  assign n15651 = ~n15597 & n15650;
  assign n15652 = n15651 ^ n15445;
  assign n15819 = n15818 ^ n15652;
  assign n15828 = n15827 ^ n15819;
  assign n15647 = n15606 ^ n15434;
  assign n15648 = n15607 & n15647;
  assign n15649 = n15648 ^ n15434;
  assign n15829 = n15828 ^ n15649;
  assign n15641 = n1746 & ~n10281;
  assign n15642 = x127 & n1750;
  assign n15643 = x126 & n1871;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = ~n15641 & n15644;
  assign n15646 = n15645 ^ x23;
  assign n15830 = n15829 ^ n15646;
  assign n15638 = n15608 ^ n15431;
  assign n15639 = ~n15617 & n15638;
  assign n15640 = n15639 ^ n15616;
  assign n15831 = n15830 ^ n15640;
  assign n15842 = n15841 ^ n15831;
  assign n16030 = n2102 & ~n10570;
  assign n16031 = x124 & n2112;
  assign n16032 = x125 & n2105;
  assign n16033 = ~n16031 & ~n16032;
  assign n16034 = x126 & n2381;
  assign n16035 = n16033 & ~n16034;
  assign n16036 = ~n16030 & n16035;
  assign n16037 = n16036 ^ x26;
  assign n16020 = n2527 & n9691;
  assign n16021 = x121 & n2690;
  assign n16022 = x123 & n2693;
  assign n16023 = ~n16021 & ~n16022;
  assign n16024 = x122 & n2530;
  assign n16025 = n16023 & ~n16024;
  assign n16026 = ~n16020 & n16025;
  assign n16027 = n16026 ^ x29;
  assign n16010 = n3009 & n8820;
  assign n16011 = x118 & n3181;
  assign n16012 = x119 & n3013;
  assign n16013 = ~n16011 & ~n16012;
  assign n16014 = x120 & n3183;
  assign n16015 = n16013 & ~n16014;
  assign n16016 = ~n16010 & n16015;
  assign n16017 = n16016 ^ x32;
  assign n16000 = n3522 & n7987;
  assign n16001 = x115 & n3699;
  assign n16002 = x116 & n3526;
  assign n16003 = ~n16001 & ~n16002;
  assign n16004 = x117 & n3701;
  assign n16005 = n16003 & ~n16004;
  assign n16006 = ~n16000 & n16005;
  assign n16007 = n16006 ^ x35;
  assign n15990 = n4040 & n7220;
  assign n15991 = x112 & n4267;
  assign n15992 = x113 & n4044;
  assign n15993 = ~n15991 & ~n15992;
  assign n15994 = x114 & n4270;
  assign n15995 = n15993 & ~n15994;
  assign n15996 = ~n15990 & n15995;
  assign n15997 = n15996 ^ x38;
  assign n15980 = n4643 & n6478;
  assign n15981 = x109 & n4653;
  assign n15982 = x111 & n5046;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = x110 & n4646;
  assign n15985 = n15983 & ~n15984;
  assign n15986 = ~n15980 & n15985;
  assign n15987 = n15986 ^ x41;
  assign n15967 = n5117 & n5942;
  assign n15968 = x103 & n6186;
  assign n15969 = x105 & n6406;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = x104 & n5947;
  assign n15972 = n15970 & ~n15971;
  assign n15973 = ~n15967 & n15972;
  assign n15974 = n15973 ^ x47;
  assign n15964 = n15743 ^ n15681;
  assign n15965 = ~n15752 & n15964;
  assign n15966 = n15965 ^ n15751;
  assign n15975 = n15974 ^ n15966;
  assign n15954 = n4509 & n6626;
  assign n15955 = x100 & n6884;
  assign n15956 = x102 & n6888;
  assign n15957 = ~n15955 & ~n15956;
  assign n15958 = x101 & n6630;
  assign n15959 = n15957 & ~n15958;
  assign n15960 = ~n15954 & n15959;
  assign n15961 = n15960 ^ x50;
  assign n15951 = n15733 ^ n15684;
  assign n15952 = ~n15742 & n15951;
  assign n15953 = n15952 ^ n15741;
  assign n15962 = n15961 ^ n15953;
  assign n15941 = n3943 & n7395;
  assign n15942 = x97 & n7650;
  assign n15943 = x98 & n7400;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = x99 & n7652;
  assign n15946 = n15944 & ~n15945;
  assign n15947 = ~n15941 & n15946;
  assign n15948 = n15947 ^ x53;
  assign n15938 = n15723 ^ n15687;
  assign n15939 = ~n15732 & n15938;
  assign n15940 = n15939 ^ n15731;
  assign n15949 = n15948 ^ n15940;
  assign n15928 = n3403 & n8171;
  assign n15929 = x94 & n8181;
  assign n15930 = x96 & n8732;
  assign n15931 = ~n15929 & ~n15930;
  assign n15932 = x95 & n8174;
  assign n15933 = n15931 & ~n15932;
  assign n15934 = ~n15928 & n15933;
  assign n15935 = n15934 ^ x56;
  assign n15925 = n15713 ^ n15690;
  assign n15926 = n15722 & n15925;
  assign n15927 = n15926 ^ n15721;
  assign n15936 = n15935 ^ n15927;
  assign n15915 = n2901 & n9002;
  assign n15916 = x91 & n9012;
  assign n15917 = x92 & n9005;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = x93 & n9557;
  assign n15920 = n15918 & ~n15919;
  assign n15921 = ~n15915 & n15920;
  assign n15922 = n15921 ^ x59;
  assign n15912 = n15703 ^ n15693;
  assign n15913 = ~n15712 & ~n15912;
  assign n15914 = n15913 ^ n15711;
  assign n15923 = n15922 ^ n15914;
  assign n15903 = n2448 & n9878;
  assign n15904 = x88 & n9888;
  assign n15905 = x89 & n9881;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = x90 & n10501;
  assign n15908 = n15906 & ~n15907;
  assign n15909 = ~n15903 & n15908;
  assign n15910 = n15909 ^ x62;
  assign n15895 = n1790 ^ x63;
  assign n15896 = n15895 ^ n1790;
  assign n15897 = n1790 ^ n1648;
  assign n15898 = n15897 ^ n1790;
  assign n15899 = n15896 & n15898;
  assign n15900 = n15899 ^ n1790;
  assign n15901 = ~n10177 & n15900;
  assign n15902 = n15901 ^ n1790;
  assign n15911 = n15910 ^ n15902;
  assign n15924 = n15923 ^ n15911;
  assign n15937 = n15936 ^ n15924;
  assign n15950 = n15949 ^ n15937;
  assign n15963 = n15962 ^ n15950;
  assign n15976 = n15975 ^ n15963;
  assign n15892 = n15756 ^ n15753;
  assign n15893 = n15765 & n15892;
  assign n15894 = n15893 ^ n15764;
  assign n15977 = n15976 ^ n15894;
  assign n15884 = n5262 & n5792;
  assign n15885 = x106 & n5488;
  assign n15886 = x107 & n5266;
  assign n15887 = ~n15885 & ~n15886;
  assign n15888 = x108 & n5491;
  assign n15889 = n15887 & ~n15888;
  assign n15890 = ~n15884 & n15889;
  assign n15891 = n15890 ^ x44;
  assign n15978 = n15977 ^ n15891;
  assign n15881 = n15775 ^ n15766;
  assign n15882 = n15767 & ~n15881;
  assign n15883 = n15882 ^ n15775;
  assign n15979 = n15978 ^ n15883;
  assign n15988 = n15987 ^ n15979;
  assign n15878 = n15784 ^ n15675;
  assign n15879 = n15785 & n15878;
  assign n15880 = n15879 ^ n15675;
  assign n15989 = n15988 ^ n15880;
  assign n15998 = n15997 ^ n15989;
  assign n15875 = n15795 ^ n15672;
  assign n15876 = n15787 & n15875;
  assign n15877 = n15876 ^ n15795;
  assign n15999 = n15998 ^ n15877;
  assign n16008 = n16007 ^ n15999;
  assign n15872 = n15805 ^ n15669;
  assign n15873 = n15797 & n15872;
  assign n15874 = n15873 ^ n15805;
  assign n16009 = n16008 ^ n15874;
  assign n16018 = n16017 ^ n16009;
  assign n15869 = n15806 ^ n15663;
  assign n15870 = ~n15807 & n15869;
  assign n15871 = n15870 ^ n15666;
  assign n16019 = n16018 ^ n15871;
  assign n16028 = n16027 ^ n16019;
  assign n15866 = n15817 ^ n15655;
  assign n15867 = n15809 & n15866;
  assign n15868 = n15867 ^ n15817;
  assign n16029 = n16028 ^ n15868;
  assign n16038 = n16037 ^ n16029;
  assign n15863 = n15827 ^ n15818;
  assign n15864 = n15819 & ~n15863;
  assign n15865 = n15864 ^ n15827;
  assign n16039 = n16038 ^ n15865;
  assign n15849 = x127 & n1625;
  assign n15850 = ~x23 & ~n15849;
  assign n15851 = n15850 ^ x22;
  assign n15852 = n1507 & n11409;
  assign n15853 = n15852 ^ n15850;
  assign n15854 = ~n15850 & n15853;
  assign n15855 = n15854 ^ n15850;
  assign n15856 = x127 & n1870;
  assign n15857 = ~n15855 & ~n15856;
  assign n15858 = n15857 ^ n15854;
  assign n15859 = n15858 ^ n15850;
  assign n15860 = n15859 ^ n15852;
  assign n15861 = ~n15851 & n15860;
  assign n15862 = n15861 ^ x22;
  assign n16040 = n16039 ^ n15862;
  assign n15846 = n15828 ^ n15646;
  assign n15847 = ~n15829 & n15846;
  assign n15848 = n15847 ^ n15649;
  assign n16041 = n16040 ^ n15848;
  assign n15843 = n15841 ^ n15640;
  assign n15844 = n15831 & ~n15843;
  assign n15845 = n15844 ^ n15841;
  assign n16042 = n16041 ^ n15845;
  assign n16232 = n15848 ^ n15845;
  assign n16233 = ~n16041 & ~n16232;
  assign n16234 = n16233 ^ n15845;
  assign n16221 = n2102 & ~n10855;
  assign n16222 = x125 & n2112;
  assign n16223 = x126 & n2105;
  assign n16224 = ~n16222 & ~n16223;
  assign n16225 = x127 & n2381;
  assign n16226 = n16224 & ~n16225;
  assign n16227 = ~n16221 & n16226;
  assign n16228 = n16227 ^ x26;
  assign n16211 = n2527 & n9999;
  assign n16212 = x122 & n2690;
  assign n16213 = x123 & n2530;
  assign n16214 = ~n16212 & ~n16213;
  assign n16215 = x124 & n2693;
  assign n16216 = n16214 & ~n16215;
  assign n16217 = ~n16211 & n16216;
  assign n16218 = n16217 ^ x29;
  assign n16199 = n3522 & n8265;
  assign n16200 = x116 & n3699;
  assign n16201 = x118 & n3701;
  assign n16202 = ~n16200 & ~n16201;
  assign n16203 = x117 & n3526;
  assign n16204 = n16202 & ~n16203;
  assign n16205 = ~n16199 & n16204;
  assign n16206 = n16205 ^ x35;
  assign n16189 = n4040 & n7481;
  assign n16190 = x113 & n4267;
  assign n16191 = x115 & n4270;
  assign n16192 = ~n16190 & ~n16191;
  assign n16193 = x114 & n4044;
  assign n16194 = n16192 & ~n16193;
  assign n16195 = ~n16189 & n16194;
  assign n16196 = n16195 ^ x38;
  assign n16179 = n4643 & n6728;
  assign n16180 = x110 & n4653;
  assign n16181 = x112 & n5046;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = x111 & n4646;
  assign n16184 = n16182 & ~n16183;
  assign n16185 = ~n16179 & n16184;
  assign n16186 = n16185 ^ x41;
  assign n16165 = n4718 & n6626;
  assign n16166 = x101 & n6884;
  assign n16167 = x103 & n6888;
  assign n16168 = ~n16166 & ~n16167;
  assign n16169 = x102 & n6630;
  assign n16170 = n16168 & ~n16169;
  assign n16171 = ~n16165 & n16170;
  assign n16172 = n16171 ^ x50;
  assign n16162 = n15953 ^ n15950;
  assign n16163 = n15962 & n16162;
  assign n16164 = n16163 ^ n15961;
  assign n16173 = n16172 ^ n16164;
  assign n16152 = n4141 & n7395;
  assign n16153 = x98 & n7650;
  assign n16154 = x99 & n7400;
  assign n16155 = ~n16153 & ~n16154;
  assign n16156 = x100 & n7652;
  assign n16157 = n16155 & ~n16156;
  assign n16158 = ~n16152 & n16157;
  assign n16159 = n16158 ^ x53;
  assign n16149 = n15940 ^ n15937;
  assign n16150 = n15949 & n16149;
  assign n16151 = n16150 ^ n15948;
  assign n16160 = n16159 ^ n16151;
  assign n16137 = n3078 & n9002;
  assign n16138 = x92 & n9012;
  assign n16139 = x93 & n9005;
  assign n16140 = ~n16138 & ~n16139;
  assign n16141 = x94 & n9557;
  assign n16142 = n16140 & ~n16141;
  assign n16143 = ~n16137 & n16142;
  assign n16144 = n16143 ^ x59;
  assign n16134 = n15914 ^ n15911;
  assign n16135 = n15923 & n16134;
  assign n16136 = n16135 ^ n15922;
  assign n16145 = n16144 ^ n16136;
  assign n16123 = ~n15902 & ~n15910;
  assign n16124 = n15692 ^ x87;
  assign n16125 = n16124 ^ n15692;
  assign n16126 = n15692 ^ n10177;
  assign n16127 = n16126 ^ n15692;
  assign n16128 = ~n16125 & n16127;
  assign n16129 = n16128 ^ n15692;
  assign n16130 = x86 & n16129;
  assign n16131 = n16130 ^ n15692;
  assign n16132 = ~n16123 & ~n16131;
  assign n16114 = n2607 & n9878;
  assign n16115 = x89 & n9888;
  assign n16116 = x91 & n10501;
  assign n16117 = ~n16115 & ~n16116;
  assign n16118 = x90 & n9881;
  assign n16119 = n16117 & ~n16118;
  assign n16120 = ~n16114 & n16119;
  assign n16121 = n16120 ^ x62;
  assign n16105 = n1909 ^ x63;
  assign n16106 = n16105 ^ n1909;
  assign n16107 = n1909 ^ n1790;
  assign n16108 = n16107 ^ n1909;
  assign n16109 = n16106 & n16108;
  assign n16110 = n16109 ^ n1909;
  assign n16111 = ~n10177 & n16110;
  assign n16112 = n16111 ^ n1909;
  assign n16113 = n16112 ^ x23;
  assign n16122 = n16121 ^ n16113;
  assign n16133 = n16132 ^ n16122;
  assign n16146 = n16145 ^ n16133;
  assign n16097 = n3585 & n8171;
  assign n16098 = x95 & n8181;
  assign n16099 = x96 & n8174;
  assign n16100 = ~n16098 & ~n16099;
  assign n16101 = x97 & n8732;
  assign n16102 = n16100 & ~n16101;
  assign n16103 = ~n16097 & n16102;
  assign n16104 = n16103 ^ x56;
  assign n16147 = n16146 ^ n16104;
  assign n16094 = n15927 ^ n15924;
  assign n16095 = n15936 & n16094;
  assign n16096 = n16095 ^ n15935;
  assign n16148 = n16147 ^ n16096;
  assign n16161 = n16160 ^ n16148;
  assign n16174 = n16173 ^ n16161;
  assign n16091 = n15966 ^ n15963;
  assign n16092 = n15975 & n16091;
  assign n16093 = n16092 ^ n15974;
  assign n16175 = n16174 ^ n16093;
  assign n16083 = n5351 & n5942;
  assign n16084 = x104 & n6186;
  assign n16085 = x106 & n6406;
  assign n16086 = ~n16084 & ~n16085;
  assign n16087 = x105 & n5947;
  assign n16088 = n16086 & ~n16087;
  assign n16089 = ~n16083 & n16088;
  assign n16090 = n16089 ^ x47;
  assign n16176 = n16175 ^ n16090;
  assign n16075 = n5262 & n6026;
  assign n16076 = x107 & n5488;
  assign n16077 = x109 & n5491;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = x108 & n5266;
  assign n16080 = n16078 & ~n16079;
  assign n16081 = ~n16075 & n16080;
  assign n16082 = n16081 ^ x44;
  assign n16177 = n16176 ^ n16082;
  assign n16072 = n15976 ^ n15891;
  assign n16073 = ~n15977 & n16072;
  assign n16074 = n16073 ^ n15894;
  assign n16178 = n16177 ^ n16074;
  assign n16187 = n16186 ^ n16178;
  assign n16069 = n15987 ^ n15883;
  assign n16070 = n15979 & n16069;
  assign n16071 = n16070 ^ n15987;
  assign n16188 = n16187 ^ n16071;
  assign n16197 = n16196 ^ n16188;
  assign n16066 = n15997 ^ n15880;
  assign n16067 = n15989 & n16066;
  assign n16068 = n16067 ^ n15997;
  assign n16198 = n16197 ^ n16068;
  assign n16207 = n16206 ^ n16198;
  assign n16063 = n16007 ^ n15998;
  assign n16064 = n15999 & ~n16063;
  assign n16065 = n16064 ^ n16007;
  assign n16208 = n16207 ^ n16065;
  assign n16060 = n16017 ^ n15874;
  assign n16061 = n16009 & n16060;
  assign n16062 = n16061 ^ n16017;
  assign n16209 = n16208 ^ n16062;
  assign n16052 = n3009 & n9094;
  assign n16053 = x119 & n3181;
  assign n16054 = x120 & n3013;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = x121 & n3183;
  assign n16057 = n16055 & ~n16056;
  assign n16058 = ~n16052 & n16057;
  assign n16059 = n16058 ^ x32;
  assign n16210 = n16209 ^ n16059;
  assign n16219 = n16218 ^ n16210;
  assign n16049 = n16027 ^ n15871;
  assign n16050 = n16019 & n16049;
  assign n16051 = n16050 ^ n16027;
  assign n16220 = n16219 ^ n16051;
  assign n16229 = n16228 ^ n16220;
  assign n16046 = n16037 ^ n16028;
  assign n16047 = n16029 & ~n16046;
  assign n16048 = n16047 ^ n16037;
  assign n16230 = n16229 ^ n16048;
  assign n16043 = n16038 ^ n15862;
  assign n16044 = n16039 & n16043;
  assign n16045 = n16044 ^ n15862;
  assign n16231 = n16230 ^ n16045;
  assign n16235 = n16234 ^ n16231;
  assign n16412 = n2527 & n10303;
  assign n16413 = x123 & n2690;
  assign n16414 = x124 & n2530;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = x125 & n2693;
  assign n16417 = n16415 & ~n16416;
  assign n16418 = ~n16412 & n16417;
  assign n16419 = n16418 ^ x29;
  assign n16402 = n3009 & n9387;
  assign n16403 = x121 & n3013;
  assign n16404 = x120 & n3181;
  assign n16405 = ~n16403 & ~n16404;
  assign n16406 = x122 & n3183;
  assign n16407 = n16405 & ~n16406;
  assign n16408 = ~n16402 & n16407;
  assign n16409 = n16408 ^ x32;
  assign n16391 = n3522 & n8542;
  assign n16392 = x117 & n3699;
  assign n16393 = x118 & n3526;
  assign n16394 = ~n16392 & ~n16393;
  assign n16395 = x119 & n3701;
  assign n16396 = n16394 & ~n16395;
  assign n16397 = ~n16391 & n16396;
  assign n16398 = n16397 ^ x35;
  assign n16388 = n16196 ^ n16068;
  assign n16389 = ~n16197 & n16388;
  assign n16390 = n16389 ^ n16068;
  assign n16399 = n16398 ^ n16390;
  assign n16379 = n4040 & n7730;
  assign n16380 = x114 & n4267;
  assign n16381 = x116 & n4270;
  assign n16382 = ~n16380 & ~n16381;
  assign n16383 = x115 & n4044;
  assign n16384 = n16382 & ~n16383;
  assign n16385 = ~n16379 & n16384;
  assign n16386 = n16385 ^ x38;
  assign n16369 = n4643 & n6975;
  assign n16370 = x111 & n4653;
  assign n16371 = x113 & n5046;
  assign n16372 = ~n16370 & ~n16371;
  assign n16373 = x112 & n4646;
  assign n16374 = n16372 & ~n16373;
  assign n16375 = ~n16369 & n16374;
  assign n16376 = n16375 ^ x41;
  assign n16358 = n5262 & n6250;
  assign n16359 = x108 & n5488;
  assign n16360 = x110 & n5491;
  assign n16361 = ~n16359 & ~n16360;
  assign n16362 = x109 & n5266;
  assign n16363 = n16361 & ~n16362;
  assign n16364 = ~n16358 & n16363;
  assign n16365 = n16364 ^ x44;
  assign n16346 = n4912 & n6626;
  assign n16347 = x102 & n6884;
  assign n16348 = x103 & n6630;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = x104 & n6888;
  assign n16351 = n16349 & ~n16350;
  assign n16352 = ~n16346 & n16351;
  assign n16353 = n16352 ^ x50;
  assign n16343 = n16159 ^ n16148;
  assign n16344 = n16160 & ~n16343;
  assign n16345 = n16344 ^ n16151;
  assign n16354 = n16353 ^ n16345;
  assign n16333 = n4323 & n7395;
  assign n16334 = x99 & n7650;
  assign n16335 = x100 & n7400;
  assign n16336 = ~n16334 & ~n16335;
  assign n16337 = x101 & n7652;
  assign n16338 = n16336 & ~n16337;
  assign n16339 = ~n16333 & n16338;
  assign n16340 = n16339 ^ x53;
  assign n16330 = n16146 ^ n16096;
  assign n16331 = ~n16147 & n16330;
  assign n16332 = n16331 ^ n16096;
  assign n16341 = n16340 ^ n16332;
  assign n16320 = n3763 & n8171;
  assign n16321 = x96 & n8181;
  assign n16322 = x98 & n8732;
  assign n16323 = ~n16321 & ~n16322;
  assign n16324 = x97 & n8174;
  assign n16325 = n16323 & ~n16324;
  assign n16326 = ~n16320 & n16325;
  assign n16327 = n16326 ^ x56;
  assign n16310 = n3247 & n9002;
  assign n16311 = x93 & n9012;
  assign n16312 = x95 & n9557;
  assign n16313 = ~n16311 & ~n16312;
  assign n16314 = x94 & n9005;
  assign n16315 = n16313 & ~n16314;
  assign n16316 = ~n16310 & n16315;
  assign n16317 = n16316 ^ x59;
  assign n16301 = n2755 & n9878;
  assign n16302 = x90 & n9888;
  assign n16303 = x91 & n9881;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = x92 & n10501;
  assign n16306 = n16304 & ~n16305;
  assign n16307 = ~n16301 & n16306;
  assign n16308 = n16307 ^ x62;
  assign n16297 = x89 & n10177;
  assign n16298 = x88 & n12123;
  assign n16299 = ~n16297 & ~n16298;
  assign n16287 = x87 ^ x23;
  assign n16288 = x88 ^ x86;
  assign n16289 = n12123 ^ x88;
  assign n16290 = n16289 ^ x88;
  assign n16291 = n16288 & n16290;
  assign n16292 = n16291 ^ x88;
  assign n16293 = n16292 ^ x87;
  assign n16294 = ~n16287 & n16293;
  assign n16295 = n16294 ^ x87;
  assign n16296 = ~n12893 & n16295;
  assign n16300 = n16299 ^ n16296;
  assign n16309 = n16308 ^ n16300;
  assign n16318 = n16317 ^ n16309;
  assign n16284 = n16132 ^ n16121;
  assign n16285 = ~n16122 & n16284;
  assign n16286 = n16285 ^ n16132;
  assign n16319 = n16318 ^ n16286;
  assign n16328 = n16327 ^ n16319;
  assign n16281 = n16144 ^ n16133;
  assign n16282 = n16145 & ~n16281;
  assign n16283 = n16282 ^ n16136;
  assign n16329 = n16328 ^ n16283;
  assign n16342 = n16341 ^ n16329;
  assign n16355 = n16354 ^ n16342;
  assign n16278 = n16172 ^ n16161;
  assign n16279 = n16173 & ~n16278;
  assign n16280 = n16279 ^ n16164;
  assign n16356 = n16355 ^ n16280;
  assign n16270 = n5578 & n5942;
  assign n16271 = x105 & n6186;
  assign n16272 = x107 & n6406;
  assign n16273 = ~n16271 & ~n16272;
  assign n16274 = x106 & n5947;
  assign n16275 = n16273 & ~n16274;
  assign n16276 = ~n16270 & n16275;
  assign n16277 = n16276 ^ x47;
  assign n16357 = n16356 ^ n16277;
  assign n16366 = n16365 ^ n16357;
  assign n16267 = n16174 ^ n16090;
  assign n16268 = n16175 & ~n16267;
  assign n16269 = n16268 ^ n16093;
  assign n16367 = n16366 ^ n16269;
  assign n16264 = n16082 ^ n16074;
  assign n16265 = n16177 & ~n16264;
  assign n16266 = n16265 ^ n16176;
  assign n16368 = n16367 ^ n16266;
  assign n16377 = n16376 ^ n16368;
  assign n16261 = n16178 ^ n16071;
  assign n16262 = n16187 & ~n16261;
  assign n16263 = n16262 ^ n16186;
  assign n16378 = n16377 ^ n16263;
  assign n16387 = n16386 ^ n16378;
  assign n16400 = n16399 ^ n16387;
  assign n16258 = n16206 ^ n16065;
  assign n16259 = ~n16207 & n16258;
  assign n16260 = n16259 ^ n16065;
  assign n16401 = n16400 ^ n16260;
  assign n16410 = n16409 ^ n16401;
  assign n16255 = n16208 ^ n16059;
  assign n16256 = n16209 & ~n16255;
  assign n16257 = n16256 ^ n16062;
  assign n16411 = n16410 ^ n16257;
  assign n16420 = n16419 ^ n16411;
  assign n16252 = n16218 ^ n16051;
  assign n16253 = ~n16219 & n16252;
  assign n16254 = n16253 ^ n16051;
  assign n16421 = n16420 ^ n16254;
  assign n16246 = n2102 & ~n10281;
  assign n16247 = x127 & n2105;
  assign n16248 = x126 & n2112;
  assign n16249 = ~n16247 & ~n16248;
  assign n16250 = ~n16246 & n16249;
  assign n16251 = n16250 ^ x26;
  assign n16422 = n16421 ^ n16251;
  assign n16240 = n16220 ^ n16048;
  assign n16241 = n16048 ^ n16045;
  assign n16242 = ~n16240 & n16241;
  assign n16236 = ~n16045 & n16048;
  assign n16237 = n16220 & n16228;
  assign n16238 = ~n16236 & ~n16237;
  assign n16239 = n16238 ^ n16234;
  assign n16243 = n16242 ^ n16239;
  assign n16244 = n16231 & ~n16243;
  assign n16245 = n16244 ^ n16239;
  assign n16423 = n16422 ^ n16245;
  assign n16609 = ~n16048 & ~n16228;
  assign n16610 = n16422 & ~n16609;
  assign n16611 = n16220 ^ n16045;
  assign n16612 = n16234 ^ n16220;
  assign n16613 = ~n16611 & n16612;
  assign n16614 = n16613 ^ n16045;
  assign n16615 = ~n16610 & n16614;
  assign n16616 = n16048 & n16228;
  assign n16617 = n16045 & ~n16220;
  assign n16618 = n16422 & ~n16617;
  assign n16619 = ~n16616 & ~n16618;
  assign n16620 = n16234 & n16619;
  assign n16621 = n16228 ^ n16048;
  assign n16622 = ~n16045 & n16220;
  assign n16623 = n16622 ^ n16048;
  assign n16624 = n16621 & n16623;
  assign n16625 = n16624 ^ n16048;
  assign n16626 = ~n16422 & ~n16625;
  assign n16627 = ~n16620 & ~n16626;
  assign n16628 = ~n16615 & n16627;
  assign n16597 = n2527 & ~n10570;
  assign n16598 = x124 & n2690;
  assign n16599 = x126 & n2693;
  assign n16600 = ~n16598 & ~n16599;
  assign n16601 = x125 & n2530;
  assign n16602 = n16600 & ~n16601;
  assign n16603 = ~n16597 & n16602;
  assign n16604 = n16603 ^ x29;
  assign n16587 = n3009 & n9691;
  assign n16588 = x121 & n3181;
  assign n16589 = x122 & n3013;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = x123 & n3183;
  assign n16592 = n16590 & ~n16591;
  assign n16593 = ~n16587 & n16592;
  assign n16594 = n16593 ^ x32;
  assign n16575 = n4040 & n7987;
  assign n16576 = x115 & n4267;
  assign n16577 = x117 & n4270;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = x116 & n4044;
  assign n16580 = n16578 & ~n16579;
  assign n16581 = ~n16575 & n16580;
  assign n16582 = n16581 ^ x38;
  assign n16565 = n4643 & n7220;
  assign n16566 = x112 & n4653;
  assign n16567 = x113 & n4646;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = x114 & n5046;
  assign n16570 = n16568 & ~n16569;
  assign n16571 = ~n16565 & n16570;
  assign n16572 = n16571 ^ x41;
  assign n16555 = n5262 & n6478;
  assign n16556 = x109 & n5488;
  assign n16557 = x111 & n5491;
  assign n16558 = ~n16556 & ~n16557;
  assign n16559 = x110 & n5266;
  assign n16560 = n16558 & ~n16559;
  assign n16561 = ~n16555 & n16560;
  assign n16562 = n16561 ^ x44;
  assign n16544 = n5792 & n5942;
  assign n16545 = x106 & n6186;
  assign n16546 = x107 & n5947;
  assign n16547 = ~n16545 & ~n16546;
  assign n16548 = x108 & n6406;
  assign n16549 = n16547 & ~n16548;
  assign n16550 = ~n16544 & n16549;
  assign n16551 = n16550 ^ x47;
  assign n16535 = n5117 & n6626;
  assign n16536 = x103 & n6884;
  assign n16537 = x104 & n6630;
  assign n16538 = ~n16536 & ~n16537;
  assign n16539 = x105 & n6888;
  assign n16540 = n16538 & ~n16539;
  assign n16541 = ~n16535 & n16540;
  assign n16542 = n16541 ^ x50;
  assign n16524 = n4509 & n7395;
  assign n16525 = x101 & n7400;
  assign n16526 = x100 & n7650;
  assign n16527 = ~n16525 & ~n16526;
  assign n16528 = x102 & n7652;
  assign n16529 = n16527 & ~n16528;
  assign n16530 = ~n16524 & n16529;
  assign n16531 = n16530 ^ x53;
  assign n16514 = n3943 & n8171;
  assign n16515 = x97 & n8181;
  assign n16516 = x99 & n8732;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = x98 & n8174;
  assign n16519 = n16517 & ~n16518;
  assign n16520 = ~n16514 & n16519;
  assign n16521 = n16520 ^ x56;
  assign n16505 = n3403 & n9002;
  assign n16506 = x94 & n9012;
  assign n16507 = x95 & n9005;
  assign n16508 = ~n16506 & ~n16507;
  assign n16509 = x96 & n9557;
  assign n16510 = n16508 & ~n16509;
  assign n16511 = ~n16505 & n16510;
  assign n16512 = n16511 ^ x59;
  assign n16495 = n2901 & n9878;
  assign n16496 = x91 & n9888;
  assign n16497 = x92 & n9881;
  assign n16498 = ~n16496 & ~n16497;
  assign n16499 = x93 & n10501;
  assign n16500 = n16498 & ~n16499;
  assign n16501 = ~n16495 & n16500;
  assign n16502 = n16501 ^ x62;
  assign n16475 = n16298 ^ x90;
  assign n16476 = n16475 ^ n16298;
  assign n16477 = n16298 ^ n10177;
  assign n16478 = n16477 ^ n16298;
  assign n16479 = ~n16476 & n16478;
  assign n16480 = n16479 ^ n16298;
  assign n16481 = x89 & n16480;
  assign n16482 = n16481 ^ n16298;
  assign n16483 = n10177 ^ x89;
  assign n16484 = n2165 ^ x90;
  assign n16485 = n16484 ^ n16483;
  assign n16486 = x88 ^ x63;
  assign n16487 = ~x88 & ~n16486;
  assign n16488 = n16487 ^ x90;
  assign n16489 = n16488 ^ x88;
  assign n16490 = n16485 & ~n16489;
  assign n16491 = n16490 ^ n16487;
  assign n16492 = n16491 ^ x88;
  assign n16493 = n16483 & ~n16492;
  assign n16494 = ~n16482 & ~n16493;
  assign n16503 = n16502 ^ n16494;
  assign n16472 = n16308 ^ n16296;
  assign n16473 = ~n16300 & ~n16472;
  assign n16474 = n16473 ^ n16308;
  assign n16504 = n16503 ^ n16474;
  assign n16513 = n16512 ^ n16504;
  assign n16522 = n16521 ^ n16513;
  assign n16469 = n16309 ^ n16286;
  assign n16470 = n16318 & ~n16469;
  assign n16471 = n16470 ^ n16317;
  assign n16523 = n16522 ^ n16471;
  assign n16532 = n16531 ^ n16523;
  assign n16466 = n16319 ^ n16283;
  assign n16467 = n16328 & ~n16466;
  assign n16468 = n16467 ^ n16327;
  assign n16533 = n16532 ^ n16468;
  assign n16463 = n16332 ^ n16329;
  assign n16464 = n16341 & ~n16463;
  assign n16465 = n16464 ^ n16340;
  assign n16534 = n16533 ^ n16465;
  assign n16543 = n16542 ^ n16534;
  assign n16552 = n16551 ^ n16543;
  assign n16460 = n16345 ^ n16342;
  assign n16461 = n16354 & ~n16460;
  assign n16462 = n16461 ^ n16353;
  assign n16553 = n16552 ^ n16462;
  assign n16457 = n16355 ^ n16277;
  assign n16458 = n16356 & ~n16457;
  assign n16459 = n16458 ^ n16280;
  assign n16554 = n16553 ^ n16459;
  assign n16563 = n16562 ^ n16554;
  assign n16454 = n16365 ^ n16269;
  assign n16455 = ~n16366 & n16454;
  assign n16456 = n16455 ^ n16269;
  assign n16564 = n16563 ^ n16456;
  assign n16573 = n16572 ^ n16564;
  assign n16451 = n16376 ^ n16266;
  assign n16452 = ~n16368 & n16451;
  assign n16453 = n16452 ^ n16376;
  assign n16574 = n16573 ^ n16453;
  assign n16583 = n16582 ^ n16574;
  assign n16448 = n16386 ^ n16263;
  assign n16449 = ~n16378 & n16448;
  assign n16450 = n16449 ^ n16386;
  assign n16584 = n16583 ^ n16450;
  assign n16440 = n3522 & n8820;
  assign n16441 = x118 & n3699;
  assign n16442 = x119 & n3526;
  assign n16443 = ~n16441 & ~n16442;
  assign n16444 = x120 & n3701;
  assign n16445 = n16443 & ~n16444;
  assign n16446 = ~n16440 & n16445;
  assign n16447 = n16446 ^ x35;
  assign n16585 = n16584 ^ n16447;
  assign n16437 = n16398 ^ n16387;
  assign n16438 = n16399 & ~n16437;
  assign n16439 = n16438 ^ n16390;
  assign n16586 = n16585 ^ n16439;
  assign n16595 = n16594 ^ n16586;
  assign n16434 = n16409 ^ n16260;
  assign n16435 = ~n16401 & n16434;
  assign n16436 = n16435 ^ n16409;
  assign n16596 = n16595 ^ n16436;
  assign n16605 = n16604 ^ n16596;
  assign n16430 = n2102 & n11409;
  assign n16431 = x127 & n2112;
  assign n16432 = ~n16430 & ~n16431;
  assign n16433 = n16432 ^ x26;
  assign n16606 = n16605 ^ n16433;
  assign n16427 = n16419 ^ n16410;
  assign n16428 = ~n16411 & n16427;
  assign n16429 = n16428 ^ n16419;
  assign n16607 = n16606 ^ n16429;
  assign n16424 = n16420 ^ n16251;
  assign n16425 = n16421 & ~n16424;
  assign n16426 = n16425 ^ n16254;
  assign n16608 = n16607 ^ n16426;
  assign n16629 = n16628 ^ n16608;
  assign n16794 = ~n16426 & ~n16429;
  assign n16795 = n16628 & ~n16794;
  assign n16796 = n16426 & n16429;
  assign n16797 = n16796 ^ n16433;
  assign n16798 = n16606 & ~n16797;
  assign n16799 = n16798 ^ n16605;
  assign n16800 = n16795 & n16799;
  assign n16801 = n16433 & n16605;
  assign n16802 = n16794 & ~n16801;
  assign n16803 = ~n16433 & ~n16605;
  assign n16804 = ~n16796 & n16803;
  assign n16805 = ~n16802 & ~n16804;
  assign n16806 = ~n16628 & ~n16805;
  assign n16807 = n16796 ^ n16794;
  assign n16808 = n16794 ^ n16433;
  assign n16809 = n16808 ^ n16794;
  assign n16810 = n16807 & n16809;
  assign n16811 = n16810 ^ n16794;
  assign n16812 = ~n16606 & n16811;
  assign n16813 = ~n16806 & ~n16812;
  assign n16814 = ~n16800 & n16813;
  assign n16784 = n2527 & ~n10855;
  assign n16785 = x125 & n2690;
  assign n16786 = x126 & n2530;
  assign n16787 = ~n16785 & ~n16786;
  assign n16788 = x127 & n2693;
  assign n16789 = n16787 & ~n16788;
  assign n16790 = ~n16784 & n16789;
  assign n16791 = n16790 ^ x29;
  assign n16774 = n3009 & n9999;
  assign n16775 = x122 & n3181;
  assign n16776 = x123 & n3013;
  assign n16777 = ~n16775 & ~n16776;
  assign n16778 = x124 & n3183;
  assign n16779 = n16777 & ~n16778;
  assign n16780 = ~n16774 & n16779;
  assign n16781 = n16780 ^ x32;
  assign n16762 = n4040 & n8265;
  assign n16763 = x116 & n4267;
  assign n16764 = x118 & n4270;
  assign n16765 = ~n16763 & ~n16764;
  assign n16766 = x117 & n4044;
  assign n16767 = n16765 & ~n16766;
  assign n16768 = ~n16762 & n16767;
  assign n16769 = n16768 ^ x38;
  assign n16752 = n4643 & n7481;
  assign n16753 = x113 & n4653;
  assign n16754 = x115 & n5046;
  assign n16755 = ~n16753 & ~n16754;
  assign n16756 = x114 & n4646;
  assign n16757 = n16755 & ~n16756;
  assign n16758 = ~n16752 & n16757;
  assign n16759 = n16758 ^ x41;
  assign n16742 = n5262 & n6728;
  assign n16743 = x110 & n5488;
  assign n16744 = x112 & n5491;
  assign n16745 = ~n16743 & ~n16744;
  assign n16746 = x111 & n5266;
  assign n16747 = n16745 & ~n16746;
  assign n16748 = ~n16742 & n16747;
  assign n16749 = n16748 ^ x44;
  assign n16730 = n5351 & n6626;
  assign n16731 = x104 & n6884;
  assign n16732 = x106 & n6888;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = x105 & n6630;
  assign n16735 = n16733 & ~n16734;
  assign n16736 = ~n16730 & n16735;
  assign n16737 = n16736 ^ x50;
  assign n16727 = n16542 ^ n16533;
  assign n16728 = ~n16534 & n16727;
  assign n16729 = n16728 ^ n16542;
  assign n16738 = n16737 ^ n16729;
  assign n16717 = n4718 & n7395;
  assign n16718 = x101 & n7650;
  assign n16719 = x103 & n7652;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = x102 & n7400;
  assign n16722 = n16720 & ~n16721;
  assign n16723 = ~n16717 & n16722;
  assign n16724 = n16723 ^ x53;
  assign n16714 = n16523 ^ n16468;
  assign n16715 = n16532 & ~n16714;
  assign n16716 = n16715 ^ n16531;
  assign n16725 = n16724 ^ n16716;
  assign n16704 = n4141 & n8171;
  assign n16705 = x98 & n8181;
  assign n16706 = x100 & n8732;
  assign n16707 = ~n16705 & ~n16706;
  assign n16708 = x99 & n8174;
  assign n16709 = n16707 & ~n16708;
  assign n16710 = ~n16704 & n16709;
  assign n16711 = n16710 ^ x56;
  assign n16694 = n3585 & n9002;
  assign n16695 = x95 & n9012;
  assign n16696 = x96 & n9005;
  assign n16697 = ~n16695 & ~n16696;
  assign n16698 = x97 & n9557;
  assign n16699 = n16697 & ~n16698;
  assign n16700 = ~n16694 & n16699;
  assign n16701 = n16700 ^ x59;
  assign n16683 = n2299 ^ x63;
  assign n16684 = n16683 ^ n2299;
  assign n16685 = n2299 ^ n2165;
  assign n16686 = n16685 ^ n2299;
  assign n16687 = n16684 & n16686;
  assign n16688 = n16687 ^ n2299;
  assign n16689 = ~n10177 & n16688;
  assign n16690 = n16689 ^ n2299;
  assign n16691 = n16690 ^ x26;
  assign n16681 = n16494 & ~n16502;
  assign n16682 = n16681 ^ n16482;
  assign n16692 = n16691 ^ n16682;
  assign n16673 = n3078 & n9878;
  assign n16674 = x92 & n9888;
  assign n16675 = x93 & n9881;
  assign n16676 = ~n16674 & ~n16675;
  assign n16677 = x94 & n10501;
  assign n16678 = n16676 & ~n16677;
  assign n16679 = ~n16673 & n16678;
  assign n16680 = n16679 ^ x62;
  assign n16693 = n16692 ^ n16680;
  assign n16702 = n16701 ^ n16693;
  assign n16670 = n16512 ^ n16474;
  assign n16671 = ~n16504 & n16670;
  assign n16672 = n16671 ^ n16512;
  assign n16703 = n16702 ^ n16672;
  assign n16712 = n16711 ^ n16703;
  assign n16667 = n16513 ^ n16471;
  assign n16668 = n16522 & ~n16667;
  assign n16669 = n16668 ^ n16521;
  assign n16713 = n16712 ^ n16669;
  assign n16726 = n16725 ^ n16713;
  assign n16739 = n16738 ^ n16726;
  assign n16659 = n5942 & n6026;
  assign n16660 = x107 & n6186;
  assign n16661 = x108 & n5947;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = x109 & n6406;
  assign n16664 = n16662 & ~n16663;
  assign n16665 = ~n16659 & n16664;
  assign n16666 = n16665 ^ x47;
  assign n16740 = n16739 ^ n16666;
  assign n16656 = n16543 ^ n16462;
  assign n16657 = n16552 & ~n16656;
  assign n16658 = n16657 ^ n16551;
  assign n16741 = n16740 ^ n16658;
  assign n16750 = n16749 ^ n16741;
  assign n16653 = n16562 ^ n16459;
  assign n16654 = ~n16554 & n16653;
  assign n16655 = n16654 ^ n16562;
  assign n16751 = n16750 ^ n16655;
  assign n16760 = n16759 ^ n16751;
  assign n16650 = n16572 ^ n16563;
  assign n16651 = ~n16564 & n16650;
  assign n16652 = n16651 ^ n16572;
  assign n16761 = n16760 ^ n16652;
  assign n16770 = n16769 ^ n16761;
  assign n16647 = n16582 ^ n16573;
  assign n16648 = ~n16574 & n16647;
  assign n16649 = n16648 ^ n16582;
  assign n16771 = n16770 ^ n16649;
  assign n16644 = n16450 ^ n16447;
  assign n16645 = n16584 & ~n16644;
  assign n16646 = n16645 ^ n16583;
  assign n16772 = n16771 ^ n16646;
  assign n16636 = n3522 & n9094;
  assign n16637 = x119 & n3699;
  assign n16638 = x120 & n3526;
  assign n16639 = ~n16637 & ~n16638;
  assign n16640 = x121 & n3701;
  assign n16641 = n16639 & ~n16640;
  assign n16642 = ~n16636 & n16641;
  assign n16643 = n16642 ^ x35;
  assign n16773 = n16772 ^ n16643;
  assign n16782 = n16781 ^ n16773;
  assign n16633 = n16594 ^ n16439;
  assign n16634 = ~n16586 & n16633;
  assign n16635 = n16634 ^ n16594;
  assign n16783 = n16782 ^ n16635;
  assign n16792 = n16791 ^ n16783;
  assign n16630 = n16604 ^ n16436;
  assign n16631 = ~n16596 & n16630;
  assign n16632 = n16631 ^ n16604;
  assign n16793 = n16792 ^ n16632;
  assign n16815 = n16814 ^ n16793;
  assign n16986 = ~n16793 & ~n16803;
  assign n16987 = ~n16796 & ~n16986;
  assign n16988 = ~n16795 & n16987;
  assign n16989 = ~n16793 & ~n16794;
  assign n16990 = ~n16801 & ~n16989;
  assign n16991 = ~n16628 & n16990;
  assign n16992 = n16793 & ~n16799;
  assign n16993 = ~n16991 & ~n16992;
  assign n16994 = ~n16988 & n16993;
  assign n16974 = n3009 & n10303;
  assign n16975 = x123 & n3181;
  assign n16976 = x124 & n3013;
  assign n16977 = ~n16975 & ~n16976;
  assign n16978 = x125 & n3183;
  assign n16979 = n16977 & ~n16978;
  assign n16980 = ~n16974 & n16979;
  assign n16981 = n16980 ^ x32;
  assign n16964 = n3522 & n9387;
  assign n16965 = x120 & n3699;
  assign n16966 = x121 & n3526;
  assign n16967 = ~n16965 & ~n16966;
  assign n16968 = x122 & n3701;
  assign n16969 = n16967 & ~n16968;
  assign n16970 = ~n16964 & n16969;
  assign n16971 = n16970 ^ x35;
  assign n16954 = n4040 & n8542;
  assign n16955 = x117 & n4267;
  assign n16956 = x119 & n4270;
  assign n16957 = ~n16955 & ~n16956;
  assign n16958 = x118 & n4044;
  assign n16959 = n16957 & ~n16958;
  assign n16960 = ~n16954 & n16959;
  assign n16961 = n16960 ^ x38;
  assign n16944 = n4643 & n7730;
  assign n16945 = x114 & n4653;
  assign n16946 = x115 & n4646;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = x116 & n5046;
  assign n16949 = n16947 & ~n16948;
  assign n16950 = ~n16944 & n16949;
  assign n16951 = n16950 ^ x41;
  assign n16927 = n4912 & n7395;
  assign n16928 = x102 & n7650;
  assign n16929 = x103 & n7400;
  assign n16930 = ~n16928 & ~n16929;
  assign n16931 = x104 & n7652;
  assign n16932 = n16930 & ~n16931;
  assign n16933 = ~n16927 & n16932;
  assign n16934 = n16933 ^ x53;
  assign n16917 = n4323 & n8171;
  assign n16918 = x99 & n8181;
  assign n16919 = x101 & n8732;
  assign n16920 = ~n16918 & ~n16919;
  assign n16921 = x100 & n8174;
  assign n16922 = n16920 & ~n16921;
  assign n16923 = ~n16917 & n16922;
  assign n16924 = n16923 ^ x56;
  assign n16914 = n16693 ^ n16672;
  assign n16915 = ~n16702 & n16914;
  assign n16916 = n16915 ^ n16701;
  assign n16925 = n16924 ^ n16916;
  assign n16904 = n3763 & n9002;
  assign n16905 = x96 & n9012;
  assign n16906 = x98 & n9557;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = x97 & n9005;
  assign n16909 = n16907 & ~n16908;
  assign n16910 = ~n16904 & n16909;
  assign n16911 = n16910 ^ x59;
  assign n16895 = n3247 & n9878;
  assign n16896 = x93 & n9888;
  assign n16897 = x94 & n9881;
  assign n16898 = ~n16896 & ~n16897;
  assign n16899 = x95 & n10501;
  assign n16900 = n16898 & ~n16899;
  assign n16901 = ~n16895 & n16900;
  assign n16902 = n16901 ^ x62;
  assign n16887 = n2437 ^ x92;
  assign n16888 = x92 ^ x63;
  assign n16889 = n16888 ^ x92;
  assign n16890 = n16887 & n16889;
  assign n16891 = n16890 ^ x92;
  assign n16892 = ~n10177 & n16891;
  assign n16893 = n16892 ^ x92;
  assign n16879 = x90 ^ x26;
  assign n16880 = x91 ^ x89;
  assign n16881 = ~n12123 & n16880;
  assign n16882 = n16881 ^ x89;
  assign n16883 = n16882 ^ x90;
  assign n16884 = ~n16879 & n16883;
  assign n16885 = n16884 ^ x90;
  assign n16886 = ~n12893 & n16885;
  assign n16894 = n16893 ^ n16886;
  assign n16903 = n16902 ^ n16894;
  assign n16912 = n16911 ^ n16903;
  assign n16876 = n16691 ^ n16680;
  assign n16877 = ~n16692 & ~n16876;
  assign n16878 = n16877 ^ n16682;
  assign n16913 = n16912 ^ n16878;
  assign n16926 = n16925 ^ n16913;
  assign n16935 = n16934 ^ n16926;
  assign n16873 = n16711 ^ n16669;
  assign n16874 = n16712 & n16873;
  assign n16875 = n16874 ^ n16669;
  assign n16936 = n16935 ^ n16875;
  assign n16870 = n16724 ^ n16713;
  assign n16871 = n16725 & n16870;
  assign n16872 = n16871 ^ n16716;
  assign n16937 = n16936 ^ n16872;
  assign n16862 = n5578 & n6626;
  assign n16863 = x105 & n6884;
  assign n16864 = x106 & n6630;
  assign n16865 = ~n16863 & ~n16864;
  assign n16866 = x107 & n6888;
  assign n16867 = n16865 & ~n16866;
  assign n16868 = ~n16862 & n16867;
  assign n16869 = n16868 ^ x50;
  assign n16938 = n16937 ^ n16869;
  assign n16859 = n16737 ^ n16726;
  assign n16860 = n16738 & n16859;
  assign n16861 = n16860 ^ n16729;
  assign n16939 = n16938 ^ n16861;
  assign n16851 = n5942 & n6250;
  assign n16852 = x108 & n6186;
  assign n16853 = x109 & n5947;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = x110 & n6406;
  assign n16856 = n16854 & ~n16855;
  assign n16857 = ~n16851 & n16856;
  assign n16858 = n16857 ^ x47;
  assign n16940 = n16939 ^ n16858;
  assign n16848 = n16666 ^ n16658;
  assign n16849 = ~n16740 & ~n16848;
  assign n16850 = n16849 ^ n16739;
  assign n16941 = n16940 ^ n16850;
  assign n16840 = n5262 & n6975;
  assign n16841 = x111 & n5488;
  assign n16842 = x113 & n5491;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = x112 & n5266;
  assign n16845 = n16843 & ~n16844;
  assign n16846 = ~n16840 & n16845;
  assign n16847 = n16846 ^ x44;
  assign n16942 = n16941 ^ n16847;
  assign n16837 = n16741 ^ n16655;
  assign n16838 = ~n16750 & n16837;
  assign n16839 = n16838 ^ n16749;
  assign n16943 = n16942 ^ n16839;
  assign n16952 = n16951 ^ n16943;
  assign n16834 = n16751 ^ n16652;
  assign n16835 = ~n16760 & n16834;
  assign n16836 = n16835 ^ n16759;
  assign n16953 = n16952 ^ n16836;
  assign n16962 = n16961 ^ n16953;
  assign n16831 = n16761 ^ n16649;
  assign n16832 = ~n16770 & n16831;
  assign n16833 = n16832 ^ n16769;
  assign n16963 = n16962 ^ n16833;
  assign n16972 = n16971 ^ n16963;
  assign n16828 = n16771 ^ n16643;
  assign n16829 = ~n16772 & n16828;
  assign n16830 = n16829 ^ n16646;
  assign n16973 = n16972 ^ n16830;
  assign n16982 = n16981 ^ n16973;
  assign n16825 = n16781 ^ n16635;
  assign n16826 = n16782 & n16825;
  assign n16827 = n16826 ^ n16635;
  assign n16983 = n16982 ^ n16827;
  assign n16819 = n2527 & ~n10281;
  assign n16820 = x127 & n2530;
  assign n16821 = x126 & n2690;
  assign n16822 = ~n16820 & ~n16821;
  assign n16823 = ~n16819 & n16822;
  assign n16824 = n16823 ^ x29;
  assign n16984 = n16983 ^ n16824;
  assign n16816 = n16791 ^ n16632;
  assign n16817 = n16792 & n16816;
  assign n16818 = n16817 ^ n16632;
  assign n16985 = n16984 ^ n16818;
  assign n16995 = n16994 ^ n16985;
  assign n17170 = n3009 & ~n10570;
  assign n17171 = x124 & n3181;
  assign n17172 = x125 & n3013;
  assign n17173 = ~n17171 & ~n17172;
  assign n17174 = x126 & n3183;
  assign n17175 = n17173 & ~n17174;
  assign n17176 = ~n17170 & n17175;
  assign n17177 = n17176 ^ x32;
  assign n17160 = n3522 & n9691;
  assign n17161 = x121 & n3699;
  assign n17162 = x123 & n3701;
  assign n17163 = ~n17161 & ~n17162;
  assign n17164 = x122 & n3526;
  assign n17165 = n17163 & ~n17164;
  assign n17166 = ~n17160 & n17165;
  assign n17167 = n17166 ^ x35;
  assign n17150 = n4040 & n8820;
  assign n17151 = x118 & n4267;
  assign n17152 = x120 & n4270;
  assign n17153 = ~n17151 & ~n17152;
  assign n17154 = x119 & n4044;
  assign n17155 = n17153 & ~n17154;
  assign n17156 = ~n17150 & n17155;
  assign n17157 = n17156 ^ x38;
  assign n17140 = n4643 & n7987;
  assign n17141 = x115 & n4653;
  assign n17142 = x117 & n5046;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = x116 & n4646;
  assign n17145 = n17143 & ~n17144;
  assign n17146 = ~n17140 & n17145;
  assign n17147 = n17146 ^ x41;
  assign n17128 = n5942 & n6478;
  assign n17129 = x109 & n6186;
  assign n17130 = x110 & n5947;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = x111 & n6406;
  assign n17133 = n17131 & ~n17132;
  assign n17134 = ~n17128 & n17133;
  assign n17135 = n17134 ^ x47;
  assign n17117 = n5792 & n6626;
  assign n17118 = x106 & n6884;
  assign n17119 = x107 & n6630;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = x108 & n6888;
  assign n17122 = n17120 & ~n17121;
  assign n17123 = ~n17117 & n17122;
  assign n17124 = n17123 ^ x50;
  assign n17114 = n16926 ^ n16875;
  assign n17115 = n16935 & ~n17114;
  assign n17116 = n17115 ^ n16934;
  assign n17125 = n17124 ^ n17116;
  assign n17104 = n5117 & n7395;
  assign n17105 = x103 & n7650;
  assign n17106 = x105 & n7652;
  assign n17107 = ~n17105 & ~n17106;
  assign n17108 = x104 & n7400;
  assign n17109 = n17107 & ~n17108;
  assign n17110 = ~n17104 & n17109;
  assign n17111 = n17110 ^ x53;
  assign n17101 = n16916 ^ n16913;
  assign n17102 = n16925 & ~n17101;
  assign n17103 = n17102 ^ n16924;
  assign n17112 = n17111 ^ n17103;
  assign n17091 = n4509 & n8171;
  assign n17092 = x100 & n8181;
  assign n17093 = x101 & n8174;
  assign n17094 = ~n17092 & ~n17093;
  assign n17095 = x102 & n8732;
  assign n17096 = n17094 & ~n17095;
  assign n17097 = ~n17091 & n17096;
  assign n17098 = n17097 ^ x56;
  assign n17088 = n16903 ^ n16878;
  assign n17089 = ~n16912 & ~n17088;
  assign n17090 = n17089 ^ n16911;
  assign n17099 = n17098 ^ n17090;
  assign n17079 = n3943 & n9002;
  assign n17080 = x97 & n9012;
  assign n17081 = x99 & n9557;
  assign n17082 = ~n17080 & ~n17081;
  assign n17083 = x98 & n9005;
  assign n17084 = n17082 & ~n17083;
  assign n17085 = ~n17079 & n17084;
  assign n17086 = n17085 ^ x59;
  assign n17056 = x92 & ~x93;
  assign n17057 = n17056 ^ x63;
  assign n17058 = n17057 ^ n17056;
  assign n17059 = x91 & ~x92;
  assign n17060 = n17059 ^ n17056;
  assign n17061 = n17060 ^ n17056;
  assign n17062 = n17058 & n17061;
  assign n17063 = n17062 ^ n17056;
  assign n17064 = ~n10177 & n17063;
  assign n17065 = n17064 ^ n17056;
  assign n17067 = ~x91 & x92;
  assign n17066 = ~x92 & x93;
  assign n17068 = n17067 ^ n17066;
  assign n17069 = n17068 ^ n17066;
  assign n17070 = n17066 ^ x63;
  assign n17071 = n17070 ^ n17066;
  assign n17072 = n17069 & n17071;
  assign n17073 = n17072 ^ n17066;
  assign n17074 = ~n10177 & n17073;
  assign n17075 = n17074 ^ n17066;
  assign n17076 = ~n17065 & ~n17075;
  assign n17053 = n16902 ^ n16886;
  assign n17054 = n16894 & ~n17053;
  assign n17055 = n17054 ^ n16902;
  assign n17077 = n17076 ^ n17055;
  assign n17045 = n3403 & n9878;
  assign n17046 = x94 & n9888;
  assign n17047 = x96 & n10501;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = x95 & n9881;
  assign n17050 = n17048 & ~n17049;
  assign n17051 = ~n17045 & n17050;
  assign n17052 = n17051 ^ x62;
  assign n17078 = n17077 ^ n17052;
  assign n17087 = n17086 ^ n17078;
  assign n17100 = n17099 ^ n17087;
  assign n17113 = n17112 ^ n17100;
  assign n17126 = n17125 ^ n17113;
  assign n17042 = n16936 ^ n16869;
  assign n17043 = n16937 & ~n17042;
  assign n17044 = n17043 ^ n16872;
  assign n17127 = n17126 ^ n17044;
  assign n17136 = n17135 ^ n17127;
  assign n17039 = n16938 ^ n16858;
  assign n17040 = n16939 & ~n17039;
  assign n17041 = n17040 ^ n16861;
  assign n17137 = n17136 ^ n17041;
  assign n17031 = n5262 & n7220;
  assign n17032 = x112 & n5488;
  assign n17033 = x114 & n5491;
  assign n17034 = ~n17032 & ~n17033;
  assign n17035 = x113 & n5266;
  assign n17036 = n17034 & ~n17035;
  assign n17037 = ~n17031 & n17036;
  assign n17038 = n17037 ^ x44;
  assign n17138 = n17137 ^ n17038;
  assign n17028 = n16940 ^ n16847;
  assign n17029 = ~n16941 & ~n17028;
  assign n17030 = n17029 ^ n16850;
  assign n17139 = n17138 ^ n17030;
  assign n17148 = n17147 ^ n17139;
  assign n17025 = n16951 ^ n16839;
  assign n17026 = n16943 & n17025;
  assign n17027 = n17026 ^ n16951;
  assign n17149 = n17148 ^ n17027;
  assign n17158 = n17157 ^ n17149;
  assign n17022 = n16961 ^ n16836;
  assign n17023 = n16953 & n17022;
  assign n17024 = n17023 ^ n16961;
  assign n17159 = n17158 ^ n17024;
  assign n17168 = n17167 ^ n17159;
  assign n17019 = n16971 ^ n16833;
  assign n17020 = n16963 & n17019;
  assign n17021 = n17020 ^ n16971;
  assign n17169 = n17168 ^ n17021;
  assign n17178 = n17177 ^ n17169;
  assign n17016 = n16981 ^ n16972;
  assign n17017 = n16973 & ~n17016;
  assign n17018 = n17017 ^ n16981;
  assign n17179 = n17178 ^ n17018;
  assign n17002 = x127 & n2390;
  assign n17003 = ~x29 & ~n17002;
  assign n17004 = n17003 ^ x28;
  assign n17005 = n2254 & n11409;
  assign n17006 = n17005 ^ n17003;
  assign n17007 = ~n17003 & n17006;
  assign n17008 = n17007 ^ n17003;
  assign n17009 = x127 & n2689;
  assign n17010 = ~n17008 & ~n17009;
  assign n17011 = n17010 ^ n17007;
  assign n17012 = n17011 ^ n17003;
  assign n17013 = n17012 ^ n17005;
  assign n17014 = ~n17004 & n17013;
  assign n17015 = n17014 ^ x28;
  assign n17180 = n17179 ^ n17015;
  assign n16999 = n16982 ^ n16824;
  assign n17000 = ~n16983 & n16999;
  assign n17001 = n17000 ^ n16827;
  assign n17181 = n17180 ^ n17001;
  assign n16996 = n16994 ^ n16818;
  assign n16997 = n16985 & n16996;
  assign n16998 = n16997 ^ n16994;
  assign n17182 = n17181 ^ n16998;
  assign n17336 = n17178 ^ n17015;
  assign n17337 = n17179 & n17336;
  assign n17338 = n17337 ^ n17015;
  assign n17333 = n17177 ^ n17168;
  assign n17334 = n17169 & ~n17333;
  assign n17335 = n17334 ^ n17177;
  assign n17339 = n17338 ^ n17335;
  assign n17324 = n3009 & ~n10855;
  assign n17325 = x125 & n3181;
  assign n17326 = x126 & n3013;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = x127 & n3183;
  assign n17329 = n17327 & ~n17328;
  assign n17330 = ~n17324 & n17329;
  assign n17331 = n17330 ^ x32;
  assign n17314 = n3522 & n9999;
  assign n17315 = x122 & n3699;
  assign n17316 = x124 & n3701;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = x123 & n3526;
  assign n17319 = n17317 & ~n17318;
  assign n17320 = ~n17314 & n17319;
  assign n17321 = n17320 ^ x35;
  assign n17302 = n4643 & n8265;
  assign n17303 = x116 & n4653;
  assign n17304 = x118 & n5046;
  assign n17305 = ~n17303 & ~n17304;
  assign n17306 = x117 & n4646;
  assign n17307 = n17305 & ~n17306;
  assign n17308 = ~n17302 & n17307;
  assign n17309 = n17308 ^ x41;
  assign n17292 = n5262 & n7481;
  assign n17293 = x113 & n5488;
  assign n17294 = x115 & n5491;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = x114 & n5266;
  assign n17297 = n17295 & ~n17296;
  assign n17298 = ~n17292 & n17297;
  assign n17299 = n17298 ^ x44;
  assign n17282 = n5942 & n6728;
  assign n17283 = x110 & n6186;
  assign n17284 = x111 & n5947;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = x112 & n6406;
  assign n17287 = n17285 & ~n17286;
  assign n17288 = ~n17282 & n17287;
  assign n17289 = n17288 ^ x47;
  assign n17272 = n6026 & n6626;
  assign n17273 = x107 & n6884;
  assign n17274 = x108 & n6630;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = x109 & n6888;
  assign n17277 = n17275 & ~n17276;
  assign n17278 = ~n17272 & n17277;
  assign n17279 = n17278 ^ x50;
  assign n17269 = n17116 ^ n17113;
  assign n17270 = n17125 & ~n17269;
  assign n17271 = n17270 ^ n17124;
  assign n17280 = n17279 ^ n17271;
  assign n17259 = n5351 & n7395;
  assign n17260 = x104 & n7650;
  assign n17261 = x105 & n7400;
  assign n17262 = ~n17260 & ~n17261;
  assign n17263 = x106 & n7652;
  assign n17264 = n17262 & ~n17263;
  assign n17265 = ~n17259 & n17264;
  assign n17266 = n17265 ^ x53;
  assign n17256 = n17103 ^ n17100;
  assign n17257 = n17112 & ~n17256;
  assign n17258 = n17257 ^ n17111;
  assign n17267 = n17266 ^ n17258;
  assign n17246 = n4718 & n8171;
  assign n17247 = x101 & n8181;
  assign n17248 = x103 & n8732;
  assign n17249 = ~n17247 & ~n17248;
  assign n17250 = x102 & n8174;
  assign n17251 = n17249 & ~n17250;
  assign n17252 = ~n17246 & n17251;
  assign n17253 = n17252 ^ x56;
  assign n17243 = n17090 ^ n17087;
  assign n17244 = n17099 & ~n17243;
  assign n17245 = n17244 ^ n17098;
  assign n17254 = n17253 ^ n17245;
  assign n17233 = n4141 & n9002;
  assign n17234 = x98 & n9012;
  assign n17235 = x99 & n9005;
  assign n17236 = ~n17234 & ~n17235;
  assign n17237 = x100 & n9557;
  assign n17238 = n17236 & ~n17237;
  assign n17239 = ~n17233 & n17238;
  assign n17240 = n17239 ^ x59;
  assign n17230 = n17086 ^ n17077;
  assign n17231 = ~n17078 & n17230;
  assign n17232 = n17231 ^ n17086;
  assign n17241 = n17240 ^ n17232;
  assign n17220 = n3585 & n9878;
  assign n17221 = x95 & n9888;
  assign n17222 = x96 & n9881;
  assign n17223 = ~n17221 & ~n17222;
  assign n17224 = x97 & n10501;
  assign n17225 = n17223 & ~n17224;
  assign n17226 = ~n17220 & n17225;
  assign n17227 = n17226 ^ x62;
  assign n17211 = n2744 ^ x63;
  assign n17212 = n17211 ^ n2744;
  assign n17213 = n2744 ^ n2585;
  assign n17214 = n17213 ^ n2744;
  assign n17215 = n17212 & n17214;
  assign n17216 = n17215 ^ n2744;
  assign n17217 = ~n10177 & n17216;
  assign n17218 = n17217 ^ n2744;
  assign n17219 = n17218 ^ x29;
  assign n17228 = n17227 ^ n17219;
  assign n17209 = n17055 & n17076;
  assign n17210 = n17209 ^ n17075;
  assign n17229 = n17228 ^ n17210;
  assign n17242 = n17241 ^ n17229;
  assign n17255 = n17254 ^ n17242;
  assign n17268 = n17267 ^ n17255;
  assign n17281 = n17280 ^ n17268;
  assign n17290 = n17289 ^ n17281;
  assign n17206 = n17135 ^ n17044;
  assign n17207 = ~n17127 & n17206;
  assign n17208 = n17207 ^ n17135;
  assign n17291 = n17290 ^ n17208;
  assign n17300 = n17299 ^ n17291;
  assign n17203 = n17136 ^ n17038;
  assign n17204 = n17137 & ~n17203;
  assign n17205 = n17204 ^ n17041;
  assign n17301 = n17300 ^ n17205;
  assign n17310 = n17309 ^ n17301;
  assign n17200 = n17147 ^ n17138;
  assign n17201 = n17139 & n17200;
  assign n17202 = n17201 ^ n17147;
  assign n17311 = n17310 ^ n17202;
  assign n17197 = n17157 ^ n17148;
  assign n17198 = n17149 & ~n17197;
  assign n17199 = n17198 ^ n17157;
  assign n17312 = n17311 ^ n17199;
  assign n17189 = n4040 & n9094;
  assign n17190 = x119 & n4267;
  assign n17191 = x121 & n4270;
  assign n17192 = ~n17190 & ~n17191;
  assign n17193 = x120 & n4044;
  assign n17194 = n17192 & ~n17193;
  assign n17195 = ~n17189 & n17194;
  assign n17196 = n17195 ^ x38;
  assign n17313 = n17312 ^ n17196;
  assign n17322 = n17321 ^ n17313;
  assign n17186 = n17167 ^ n17024;
  assign n17187 = n17159 & n17186;
  assign n17188 = n17187 ^ n17167;
  assign n17323 = n17322 ^ n17188;
  assign n17332 = n17331 ^ n17323;
  assign n17340 = n17339 ^ n17332;
  assign n17183 = n17001 ^ n16998;
  assign n17184 = ~n17181 & n17183;
  assign n17185 = n17184 ^ n16998;
  assign n17341 = n17340 ^ n17185;
  assign n17493 = ~n17323 & ~n17331;
  assign n17494 = ~n17335 & n17493;
  assign n17495 = n17323 & n17331;
  assign n17496 = n17335 & n17495;
  assign n17497 = ~n17494 & ~n17496;
  assign n17498 = n17339 & ~n17497;
  assign n17499 = n17335 ^ n17331;
  assign n17500 = ~n17332 & n17499;
  assign n17501 = n17500 ^ n17335;
  assign n17504 = n17338 & ~n17501;
  assign n17505 = ~n17494 & ~n17504;
  assign n17502 = ~n17338 & n17501;
  assign n17503 = ~n17496 & ~n17502;
  assign n17506 = n17505 ^ n17503;
  assign n17507 = n17185 & n17506;
  assign n17508 = n17507 ^ n17505;
  assign n17509 = ~n17498 & n17508;
  assign n17482 = n3522 & n10303;
  assign n17483 = x123 & n3699;
  assign n17484 = x125 & n3701;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = x124 & n3526;
  assign n17487 = n17485 & ~n17486;
  assign n17488 = ~n17482 & n17487;
  assign n17489 = n17488 ^ x35;
  assign n17472 = n4040 & n9387;
  assign n17473 = x120 & n4267;
  assign n17474 = x122 & n4270;
  assign n17475 = ~n17473 & ~n17474;
  assign n17476 = x121 & n4044;
  assign n17477 = n17475 & ~n17476;
  assign n17478 = ~n17472 & n17477;
  assign n17479 = n17478 ^ x38;
  assign n17460 = n5262 & n7730;
  assign n17461 = x114 & n5488;
  assign n17462 = x116 & n5491;
  assign n17463 = ~n17461 & ~n17462;
  assign n17464 = x115 & n5266;
  assign n17465 = n17463 & ~n17464;
  assign n17466 = ~n17460 & n17465;
  assign n17467 = n17466 ^ x44;
  assign n17450 = n5942 & n6975;
  assign n17451 = x111 & n6186;
  assign n17452 = x113 & n6406;
  assign n17453 = ~n17451 & ~n17452;
  assign n17454 = x112 & n5947;
  assign n17455 = n17453 & ~n17454;
  assign n17456 = ~n17450 & n17455;
  assign n17457 = n17456 ^ x47;
  assign n17439 = n6250 & n6626;
  assign n17440 = x108 & n6884;
  assign n17441 = x109 & n6630;
  assign n17442 = ~n17440 & ~n17441;
  assign n17443 = x110 & n6888;
  assign n17444 = n17442 & ~n17443;
  assign n17445 = ~n17439 & n17444;
  assign n17446 = n17445 ^ x50;
  assign n17436 = n17266 ^ n17255;
  assign n17437 = n17267 & ~n17436;
  assign n17438 = n17437 ^ n17258;
  assign n17447 = n17446 ^ n17438;
  assign n17426 = n5578 & n7395;
  assign n17427 = x106 & n7400;
  assign n17428 = x105 & n7650;
  assign n17429 = ~n17427 & ~n17428;
  assign n17430 = x107 & n7652;
  assign n17431 = n17429 & ~n17430;
  assign n17432 = ~n17426 & n17431;
  assign n17433 = n17432 ^ x53;
  assign n17423 = n17253 ^ n17242;
  assign n17424 = n17254 & ~n17423;
  assign n17425 = n17424 ^ n17245;
  assign n17434 = n17433 ^ n17425;
  assign n17413 = n4912 & n8171;
  assign n17414 = x103 & n8174;
  assign n17415 = x102 & n8181;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = x104 & n8732;
  assign n17418 = n17416 & ~n17417;
  assign n17419 = ~n17413 & n17418;
  assign n17420 = n17419 ^ x56;
  assign n17403 = n4323 & n9002;
  assign n17404 = x99 & n9012;
  assign n17405 = x101 & n9557;
  assign n17406 = ~n17404 & ~n17405;
  assign n17407 = x100 & n9005;
  assign n17408 = n17406 & ~n17407;
  assign n17409 = ~n17403 & n17408;
  assign n17410 = n17409 ^ x59;
  assign n17393 = n3763 & n9878;
  assign n17394 = x97 & n9881;
  assign n17395 = x96 & n9888;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = x98 & n10501;
  assign n17398 = n17396 & ~n17397;
  assign n17399 = ~n17393 & n17398;
  assign n17400 = n17399 ^ x62;
  assign n17383 = x93 ^ x29;
  assign n17384 = x94 ^ x92;
  assign n17385 = n12123 ^ x94;
  assign n17386 = n17385 ^ x94;
  assign n17387 = n17384 & n17386;
  assign n17388 = n17387 ^ x94;
  assign n17389 = n17388 ^ x93;
  assign n17390 = ~n17383 & n17389;
  assign n17391 = n17390 ^ x93;
  assign n17392 = ~n12893 & n17391;
  assign n17401 = n17400 ^ n17392;
  assign n17380 = x94 & n12123;
  assign n17381 = x95 & n10177;
  assign n17382 = ~n17380 & ~n17381;
  assign n17402 = n17401 ^ n17382;
  assign n17411 = n17410 ^ n17402;
  assign n17377 = n17227 ^ n17210;
  assign n17378 = ~n17228 & n17377;
  assign n17379 = n17378 ^ n17210;
  assign n17412 = n17411 ^ n17379;
  assign n17421 = n17420 ^ n17412;
  assign n17374 = n17240 ^ n17229;
  assign n17375 = n17241 & ~n17374;
  assign n17376 = n17375 ^ n17232;
  assign n17422 = n17421 ^ n17376;
  assign n17435 = n17434 ^ n17422;
  assign n17448 = n17447 ^ n17435;
  assign n17371 = n17279 ^ n17268;
  assign n17372 = n17280 & ~n17371;
  assign n17373 = n17372 ^ n17271;
  assign n17449 = n17448 ^ n17373;
  assign n17458 = n17457 ^ n17449;
  assign n17368 = n17289 ^ n17208;
  assign n17369 = ~n17290 & n17368;
  assign n17370 = n17369 ^ n17208;
  assign n17459 = n17458 ^ n17370;
  assign n17468 = n17467 ^ n17459;
  assign n17365 = n17299 ^ n17205;
  assign n17366 = ~n17300 & n17365;
  assign n17367 = n17366 ^ n17205;
  assign n17469 = n17468 ^ n17367;
  assign n17357 = n4643 & n8542;
  assign n17358 = x117 & n4653;
  assign n17359 = x118 & n4646;
  assign n17360 = ~n17358 & ~n17359;
  assign n17361 = x119 & n5046;
  assign n17362 = n17360 & ~n17361;
  assign n17363 = ~n17357 & n17362;
  assign n17364 = n17363 ^ x41;
  assign n17470 = n17469 ^ n17364;
  assign n17354 = n17309 ^ n17202;
  assign n17355 = ~n17310 & n17354;
  assign n17356 = n17355 ^ n17202;
  assign n17471 = n17470 ^ n17356;
  assign n17480 = n17479 ^ n17471;
  assign n17351 = n17311 ^ n17196;
  assign n17352 = n17312 & ~n17351;
  assign n17353 = n17352 ^ n17199;
  assign n17481 = n17480 ^ n17353;
  assign n17490 = n17489 ^ n17481;
  assign n17348 = n17321 ^ n17188;
  assign n17349 = ~n17322 & n17348;
  assign n17350 = n17349 ^ n17188;
  assign n17491 = n17490 ^ n17350;
  assign n17342 = n3009 & ~n10281;
  assign n17343 = x127 & n3013;
  assign n17344 = x126 & n3181;
  assign n17345 = ~n17343 & ~n17344;
  assign n17346 = ~n17342 & n17345;
  assign n17347 = n17346 ^ x32;
  assign n17492 = n17491 ^ n17347;
  assign n17510 = n17509 ^ n17492;
  assign n17666 = ~n17335 & n17338;
  assign n17667 = n17492 & ~n17666;
  assign n17668 = ~n17495 & ~n17667;
  assign n17669 = n17335 & ~n17338;
  assign n17670 = n17492 & ~n17493;
  assign n17671 = ~n17669 & ~n17670;
  assign n17672 = ~n17668 & ~n17671;
  assign n17673 = ~n17185 & ~n17672;
  assign n17674 = n17493 ^ n17492;
  assign n17675 = n17666 ^ n17492;
  assign n17676 = n17675 ^ n17666;
  assign n17677 = n17495 ^ n17335;
  assign n17678 = ~n17339 & n17677;
  assign n17679 = n17678 ^ n17335;
  assign n17680 = n17679 ^ n17666;
  assign n17681 = ~n17676 & n17680;
  assign n17682 = n17681 ^ n17666;
  assign n17683 = ~n17674 & ~n17682;
  assign n17684 = n17683 ^ n17493;
  assign n17685 = ~n17673 & ~n17684;
  assign n17651 = n10278 ^ x32;
  assign n17652 = n17651 ^ x32;
  assign n17653 = ~x31 & x127;
  assign n17654 = n17653 ^ x32;
  assign n17655 = ~n17652 & ~n17654;
  assign n17656 = n17655 ^ x32;
  assign n17657 = ~n2830 & ~n17656;
  assign n17658 = n3004 ^ x31;
  assign n17659 = n3008 & n17658;
  assign n17660 = x127 & n17659;
  assign n17661 = n17660 ^ x32;
  assign n17662 = ~n17657 & n17661;
  assign n17642 = n3522 & ~n10570;
  assign n17643 = x124 & n3699;
  assign n17644 = x126 & n3701;
  assign n17645 = ~n17643 & ~n17644;
  assign n17646 = x125 & n3526;
  assign n17647 = n17645 & ~n17646;
  assign n17648 = ~n17642 & n17647;
  assign n17649 = n17648 ^ x35;
  assign n17632 = n4040 & n9691;
  assign n17633 = x121 & n4267;
  assign n17634 = x122 & n4044;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = x123 & n4270;
  assign n17637 = n17635 & ~n17636;
  assign n17638 = ~n17632 & n17637;
  assign n17639 = n17638 ^ x38;
  assign n17622 = n4643 & n8820;
  assign n17623 = x118 & n4653;
  assign n17624 = x120 & n5046;
  assign n17625 = ~n17623 & ~n17624;
  assign n17626 = x119 & n4646;
  assign n17627 = n17625 & ~n17626;
  assign n17628 = ~n17622 & n17627;
  assign n17629 = n17628 ^ x41;
  assign n17612 = n5262 & n7987;
  assign n17613 = x115 & n5488;
  assign n17614 = x117 & n5491;
  assign n17615 = ~n17613 & ~n17614;
  assign n17616 = x116 & n5266;
  assign n17617 = n17615 & ~n17616;
  assign n17618 = ~n17612 & n17617;
  assign n17619 = n17618 ^ x44;
  assign n17602 = n5942 & n7220;
  assign n17603 = x112 & n6186;
  assign n17604 = x114 & n6406;
  assign n17605 = ~n17603 & ~n17604;
  assign n17606 = x113 & n5947;
  assign n17607 = n17605 & ~n17606;
  assign n17608 = ~n17602 & n17607;
  assign n17609 = n17608 ^ x47;
  assign n17592 = n6478 & n6626;
  assign n17593 = x109 & n6884;
  assign n17594 = x110 & n6630;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = x111 & n6888;
  assign n17597 = n17595 & ~n17596;
  assign n17598 = ~n17592 & n17597;
  assign n17599 = n17598 ^ x50;
  assign n17581 = n5792 & n7395;
  assign n17582 = x106 & n7650;
  assign n17583 = x107 & n7400;
  assign n17584 = ~n17582 & ~n17583;
  assign n17585 = x108 & n7652;
  assign n17586 = n17584 & ~n17585;
  assign n17587 = ~n17581 & n17586;
  assign n17588 = n17587 ^ x53;
  assign n17578 = n17412 ^ n17376;
  assign n17579 = n17421 & ~n17578;
  assign n17580 = n17579 ^ n17420;
  assign n17589 = n17588 ^ n17580;
  assign n17568 = n5117 & n8171;
  assign n17569 = x103 & n8181;
  assign n17570 = x105 & n8732;
  assign n17571 = ~n17569 & ~n17570;
  assign n17572 = x104 & n8174;
  assign n17573 = n17571 & ~n17572;
  assign n17574 = ~n17568 & n17573;
  assign n17575 = n17574 ^ x56;
  assign n17565 = n17402 ^ n17379;
  assign n17566 = n17411 & ~n17565;
  assign n17567 = n17566 ^ n17410;
  assign n17576 = n17575 ^ n17567;
  assign n17554 = n3059 ^ x63;
  assign n17555 = n17554 ^ n3059;
  assign n17556 = n3059 ^ n2890;
  assign n17557 = n17556 ^ n3059;
  assign n17558 = n17555 & n17557;
  assign n17559 = n17558 ^ n3059;
  assign n17560 = ~n10177 & n17559;
  assign n17561 = n17560 ^ n3059;
  assign n17551 = n17392 ^ n17382;
  assign n17552 = ~n17401 & ~n17551;
  assign n17553 = n17552 ^ n17400;
  assign n17562 = n17561 ^ n17553;
  assign n17543 = n3943 & n9878;
  assign n17544 = x98 & n9881;
  assign n17545 = x97 & n9888;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = x99 & n10501;
  assign n17548 = n17546 & ~n17547;
  assign n17549 = ~n17543 & n17548;
  assign n17550 = n17549 ^ x62;
  assign n17563 = n17562 ^ n17550;
  assign n17535 = n4509 & n9002;
  assign n17536 = x100 & n9012;
  assign n17537 = x101 & n9005;
  assign n17538 = ~n17536 & ~n17537;
  assign n17539 = x102 & n9557;
  assign n17540 = n17538 & ~n17539;
  assign n17541 = ~n17535 & n17540;
  assign n17542 = n17541 ^ x59;
  assign n17564 = n17563 ^ n17542;
  assign n17577 = n17576 ^ n17564;
  assign n17590 = n17589 ^ n17577;
  assign n17532 = n17433 ^ n17422;
  assign n17533 = n17434 & ~n17532;
  assign n17534 = n17533 ^ n17425;
  assign n17591 = n17590 ^ n17534;
  assign n17600 = n17599 ^ n17591;
  assign n17529 = n17446 ^ n17435;
  assign n17530 = n17447 & ~n17529;
  assign n17531 = n17530 ^ n17438;
  assign n17601 = n17600 ^ n17531;
  assign n17610 = n17609 ^ n17601;
  assign n17526 = n17457 ^ n17448;
  assign n17527 = ~n17449 & n17526;
  assign n17528 = n17527 ^ n17457;
  assign n17611 = n17610 ^ n17528;
  assign n17620 = n17619 ^ n17611;
  assign n17523 = n17467 ^ n17370;
  assign n17524 = ~n17459 & n17523;
  assign n17525 = n17524 ^ n17467;
  assign n17621 = n17620 ^ n17525;
  assign n17630 = n17629 ^ n17621;
  assign n17520 = n17468 ^ n17364;
  assign n17521 = n17469 & ~n17520;
  assign n17522 = n17521 ^ n17367;
  assign n17631 = n17630 ^ n17522;
  assign n17640 = n17639 ^ n17631;
  assign n17517 = n17479 ^ n17356;
  assign n17518 = ~n17471 & n17517;
  assign n17519 = n17518 ^ n17479;
  assign n17641 = n17640 ^ n17519;
  assign n17650 = n17649 ^ n17641;
  assign n17663 = n17662 ^ n17650;
  assign n17514 = n17489 ^ n17353;
  assign n17515 = ~n17481 & n17514;
  assign n17516 = n17515 ^ n17489;
  assign n17664 = n17663 ^ n17516;
  assign n17511 = n17490 ^ n17347;
  assign n17512 = n17491 & ~n17511;
  assign n17513 = n17512 ^ n17350;
  assign n17665 = n17664 ^ n17513;
  assign n17686 = n17685 ^ n17665;
  assign n17840 = n3522 & ~n10855;
  assign n17841 = x125 & n3699;
  assign n17842 = x126 & n3526;
  assign n17843 = ~n17841 & ~n17842;
  assign n17844 = x127 & n3701;
  assign n17845 = n17843 & ~n17844;
  assign n17846 = ~n17840 & n17845;
  assign n17847 = n17846 ^ x35;
  assign n17830 = n4040 & n9999;
  assign n17831 = x122 & n4267;
  assign n17832 = x123 & n4044;
  assign n17833 = ~n17831 & ~n17832;
  assign n17834 = x124 & n4270;
  assign n17835 = n17833 & ~n17834;
  assign n17836 = ~n17830 & n17835;
  assign n17837 = n17836 ^ x38;
  assign n17814 = n6626 & n6728;
  assign n17815 = x110 & n6884;
  assign n17816 = x111 & n6630;
  assign n17817 = ~n17815 & ~n17816;
  assign n17818 = x112 & n6888;
  assign n17819 = n17817 & ~n17818;
  assign n17820 = ~n17814 & n17819;
  assign n17821 = n17820 ^ x50;
  assign n17811 = n17599 ^ n17534;
  assign n17812 = n17591 & n17811;
  assign n17813 = n17812 ^ n17599;
  assign n17822 = n17821 ^ n17813;
  assign n17801 = n6026 & n7395;
  assign n17802 = x107 & n7650;
  assign n17803 = x109 & n7652;
  assign n17804 = ~n17802 & ~n17803;
  assign n17805 = x108 & n7400;
  assign n17806 = n17804 & ~n17805;
  assign n17807 = ~n17801 & n17806;
  assign n17808 = n17807 ^ x53;
  assign n17798 = n17588 ^ n17577;
  assign n17799 = n17589 & n17798;
  assign n17800 = n17799 ^ n17580;
  assign n17809 = n17808 ^ n17800;
  assign n17788 = n5351 & n8171;
  assign n17789 = x104 & n8181;
  assign n17790 = x105 & n8174;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = x106 & n8732;
  assign n17793 = n17791 & ~n17792;
  assign n17794 = ~n17788 & n17793;
  assign n17795 = n17794 ^ x56;
  assign n17785 = n17567 ^ n17564;
  assign n17786 = n17576 & n17785;
  assign n17787 = n17786 ^ n17575;
  assign n17796 = n17795 ^ n17787;
  assign n17775 = n4718 & n9002;
  assign n17776 = x101 & n9012;
  assign n17777 = x102 & n9005;
  assign n17778 = ~n17776 & ~n17777;
  assign n17779 = x103 & n9557;
  assign n17780 = n17778 & ~n17779;
  assign n17781 = ~n17775 & n17780;
  assign n17782 = n17781 ^ x59;
  assign n17772 = n17550 ^ n17542;
  assign n17773 = ~n17563 & ~n17772;
  assign n17774 = n17773 ^ n17562;
  assign n17783 = n17782 ^ n17774;
  assign n17750 = n17380 ^ x96;
  assign n17751 = n17750 ^ n17380;
  assign n17752 = n17380 ^ n10177;
  assign n17753 = n17752 ^ n17380;
  assign n17754 = ~n17751 & n17753;
  assign n17755 = n17754 ^ n17380;
  assign n17756 = x95 & n17755;
  assign n17757 = n17756 ^ n17380;
  assign n17758 = n17553 & ~n17757;
  assign n17759 = n10177 ^ x95;
  assign n17760 = n3059 ^ x96;
  assign n17761 = n17760 ^ n17759;
  assign n17762 = x94 ^ x63;
  assign n17763 = ~x94 & ~n17762;
  assign n17764 = n17763 ^ x96;
  assign n17765 = n17764 ^ x94;
  assign n17766 = n17761 & ~n17765;
  assign n17767 = n17766 ^ n17763;
  assign n17768 = n17767 ^ x94;
  assign n17769 = n17759 & ~n17768;
  assign n17770 = ~n17758 & ~n17769;
  assign n17741 = n4141 & n9878;
  assign n17742 = x98 & n9888;
  assign n17743 = x100 & n10501;
  assign n17744 = ~n17742 & ~n17743;
  assign n17745 = x99 & n9881;
  assign n17746 = n17744 & ~n17745;
  assign n17747 = ~n17741 & n17746;
  assign n17748 = n17747 ^ x62;
  assign n17732 = n3218 ^ x63;
  assign n17733 = n17732 ^ n3218;
  assign n17734 = n3218 ^ n3059;
  assign n17735 = n17734 ^ n3218;
  assign n17736 = n17733 & n17735;
  assign n17737 = n17736 ^ n3218;
  assign n17738 = ~n10177 & n17737;
  assign n17739 = n17738 ^ n3218;
  assign n17740 = n17739 ^ x32;
  assign n17749 = n17748 ^ n17740;
  assign n17771 = n17770 ^ n17749;
  assign n17784 = n17783 ^ n17771;
  assign n17797 = n17796 ^ n17784;
  assign n17810 = n17809 ^ n17797;
  assign n17823 = n17822 ^ n17810;
  assign n17724 = n5942 & n7481;
  assign n17725 = x113 & n6186;
  assign n17726 = x114 & n5947;
  assign n17727 = ~n17725 & ~n17726;
  assign n17728 = x115 & n6406;
  assign n17729 = n17727 & ~n17728;
  assign n17730 = ~n17724 & n17729;
  assign n17731 = n17730 ^ x47;
  assign n17824 = n17823 ^ n17731;
  assign n17721 = n17609 ^ n17531;
  assign n17722 = n17601 & n17721;
  assign n17723 = n17722 ^ n17609;
  assign n17825 = n17824 ^ n17723;
  assign n17718 = n17619 ^ n17610;
  assign n17719 = n17611 & ~n17718;
  assign n17720 = n17719 ^ n17619;
  assign n17826 = n17825 ^ n17720;
  assign n17710 = n5262 & n8265;
  assign n17711 = x116 & n5488;
  assign n17712 = x117 & n5266;
  assign n17713 = ~n17711 & ~n17712;
  assign n17714 = x118 & n5491;
  assign n17715 = n17713 & ~n17714;
  assign n17716 = ~n17710 & n17715;
  assign n17717 = n17716 ^ x44;
  assign n17827 = n17826 ^ n17717;
  assign n17707 = n17629 ^ n17620;
  assign n17708 = n17621 & ~n17707;
  assign n17709 = n17708 ^ n17629;
  assign n17828 = n17827 ^ n17709;
  assign n17699 = n4643 & n9094;
  assign n17700 = x119 & n4653;
  assign n17701 = x121 & n5046;
  assign n17702 = ~n17700 & ~n17701;
  assign n17703 = x120 & n4646;
  assign n17704 = n17702 & ~n17703;
  assign n17705 = ~n17699 & n17704;
  assign n17706 = n17705 ^ x41;
  assign n17829 = n17828 ^ n17706;
  assign n17838 = n17837 ^ n17829;
  assign n17696 = n17639 ^ n17522;
  assign n17697 = n17631 & n17696;
  assign n17698 = n17697 ^ n17639;
  assign n17839 = n17838 ^ n17698;
  assign n17848 = n17847 ^ n17839;
  assign n17693 = n17649 ^ n17640;
  assign n17694 = n17641 & ~n17693;
  assign n17695 = n17694 ^ n17649;
  assign n17849 = n17848 ^ n17695;
  assign n17690 = n17650 ^ n17516;
  assign n17691 = n17663 & n17690;
  assign n17692 = n17691 ^ n17662;
  assign n17850 = n17849 ^ n17692;
  assign n17687 = n17685 ^ n17513;
  assign n17688 = ~n17665 & n17687;
  assign n17689 = n17688 ^ n17685;
  assign n17851 = n17850 ^ n17689;
  assign n17986 = n3522 & ~n10281;
  assign n17987 = x127 & n3526;
  assign n17988 = x126 & n3699;
  assign n17989 = ~n17987 & ~n17988;
  assign n17990 = ~n17986 & n17989;
  assign n17991 = n17990 ^ x35;
  assign n17977 = n4040 & n10303;
  assign n17978 = x123 & n4267;
  assign n17979 = x125 & n4270;
  assign n17980 = ~n17978 & ~n17979;
  assign n17981 = x124 & n4044;
  assign n17982 = n17980 & ~n17981;
  assign n17983 = ~n17977 & n17982;
  assign n17984 = n17983 ^ x38;
  assign n17967 = n4643 & n9387;
  assign n17968 = x120 & n4653;
  assign n17969 = x121 & n4646;
  assign n17970 = ~n17968 & ~n17969;
  assign n17971 = x122 & n5046;
  assign n17972 = n17970 & ~n17971;
  assign n17973 = ~n17967 & n17972;
  assign n17974 = n17973 ^ x41;
  assign n17954 = n5942 & n7730;
  assign n17955 = x114 & n6186;
  assign n17956 = x116 & n6406;
  assign n17957 = ~n17955 & ~n17956;
  assign n17958 = x115 & n5947;
  assign n17959 = n17957 & ~n17958;
  assign n17960 = ~n17954 & n17959;
  assign n17961 = n17960 ^ x47;
  assign n17944 = n6626 & n6975;
  assign n17945 = x111 & n6884;
  assign n17946 = x112 & n6630;
  assign n17947 = ~n17945 & ~n17946;
  assign n17948 = x113 & n6888;
  assign n17949 = n17947 & ~n17948;
  assign n17950 = ~n17944 & n17949;
  assign n17951 = n17950 ^ x50;
  assign n17941 = n17808 ^ n17797;
  assign n17942 = n17809 & ~n17941;
  assign n17943 = n17942 ^ n17800;
  assign n17952 = n17951 ^ n17943;
  assign n17931 = n6250 & n7395;
  assign n17932 = x108 & n7650;
  assign n17933 = x110 & n7652;
  assign n17934 = ~n17932 & ~n17933;
  assign n17935 = x109 & n7400;
  assign n17936 = n17934 & ~n17935;
  assign n17937 = ~n17931 & n17936;
  assign n17938 = n17937 ^ x53;
  assign n17928 = n17795 ^ n17784;
  assign n17929 = n17796 & ~n17928;
  assign n17930 = n17929 ^ n17787;
  assign n17939 = n17938 ^ n17930;
  assign n17918 = n5578 & n8171;
  assign n17919 = x105 & n8181;
  assign n17920 = x106 & n8174;
  assign n17921 = ~n17919 & ~n17920;
  assign n17922 = x107 & n8732;
  assign n17923 = n17921 & ~n17922;
  assign n17924 = ~n17918 & n17923;
  assign n17925 = n17924 ^ x56;
  assign n17915 = n17774 ^ n17771;
  assign n17916 = ~n17783 & ~n17915;
  assign n17917 = n17916 ^ n17782;
  assign n17926 = n17925 ^ n17917;
  assign n17905 = n4912 & n9002;
  assign n17906 = x102 & n9012;
  assign n17907 = x104 & n9557;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = x103 & n9005;
  assign n17910 = n17908 & ~n17909;
  assign n17911 = ~n17905 & n17910;
  assign n17912 = n17911 ^ x59;
  assign n17895 = n4323 & n9878;
  assign n17896 = x99 & n9888;
  assign n17897 = x100 & n9881;
  assign n17898 = ~n17896 & ~n17897;
  assign n17899 = x101 & n10501;
  assign n17900 = n17898 & ~n17899;
  assign n17901 = ~n17895 & n17900;
  assign n17902 = n17901 ^ x62;
  assign n17887 = x96 ^ x32;
  assign n17888 = x97 ^ x95;
  assign n17889 = ~n12123 & n17888;
  assign n17890 = n17889 ^ x95;
  assign n17891 = n17890 ^ x96;
  assign n17892 = ~n17887 & n17891;
  assign n17893 = n17892 ^ x96;
  assign n17894 = ~n12893 & n17893;
  assign n17903 = n17902 ^ n17894;
  assign n17884 = x98 & n10177;
  assign n17885 = x97 & n12123;
  assign n17886 = ~n17884 & ~n17885;
  assign n17904 = n17903 ^ n17886;
  assign n17913 = n17912 ^ n17904;
  assign n17881 = n17770 ^ n17748;
  assign n17882 = ~n17749 & ~n17881;
  assign n17883 = n17882 ^ n17770;
  assign n17914 = n17913 ^ n17883;
  assign n17927 = n17926 ^ n17914;
  assign n17940 = n17939 ^ n17927;
  assign n17953 = n17952 ^ n17940;
  assign n17962 = n17961 ^ n17953;
  assign n17878 = n17821 ^ n17810;
  assign n17879 = n17822 & ~n17878;
  assign n17880 = n17879 ^ n17813;
  assign n17963 = n17962 ^ n17880;
  assign n17875 = n17731 ^ n17723;
  assign n17876 = n17824 & ~n17875;
  assign n17877 = n17876 ^ n17823;
  assign n17964 = n17963 ^ n17877;
  assign n17867 = n5262 & n8542;
  assign n17868 = x117 & n5488;
  assign n17869 = x118 & n5266;
  assign n17870 = ~n17868 & ~n17869;
  assign n17871 = x119 & n5491;
  assign n17872 = n17870 & ~n17871;
  assign n17873 = ~n17867 & n17872;
  assign n17874 = n17873 ^ x44;
  assign n17965 = n17964 ^ n17874;
  assign n17864 = n17825 ^ n17717;
  assign n17865 = n17826 & ~n17864;
  assign n17866 = n17865 ^ n17720;
  assign n17966 = n17965 ^ n17866;
  assign n17975 = n17974 ^ n17966;
  assign n17861 = n17827 ^ n17706;
  assign n17862 = n17828 & ~n17861;
  assign n17863 = n17862 ^ n17709;
  assign n17976 = n17975 ^ n17863;
  assign n17985 = n17984 ^ n17976;
  assign n17992 = n17991 ^ n17985;
  assign n17858 = n17837 ^ n17698;
  assign n17859 = ~n17838 & n17858;
  assign n17860 = n17859 ^ n17698;
  assign n17993 = n17992 ^ n17860;
  assign n17855 = n17839 ^ n17695;
  assign n17856 = n17848 & ~n17855;
  assign n17857 = n17856 ^ n17847;
  assign n17994 = n17993 ^ n17857;
  assign n17852 = n17692 ^ n17689;
  assign n17853 = n17850 & ~n17852;
  assign n17854 = n17853 ^ n17689;
  assign n17995 = n17994 ^ n17854;
  assign n18142 = n17985 & ~n17991;
  assign n18143 = n17860 ^ n17857;
  assign n18144 = ~n17985 & n17991;
  assign n18145 = n18144 ^ n17860;
  assign n18146 = n18143 & ~n18145;
  assign n18147 = n18146 ^ n17857;
  assign n18148 = ~n18142 & n18147;
  assign n18136 = n17857 & n17860;
  assign n18137 = ~n17857 & ~n17860;
  assign n18138 = n18137 ^ n17985;
  assign n18139 = ~n17992 & ~n18138;
  assign n18140 = n18139 ^ n17991;
  assign n18141 = ~n18136 & ~n18140;
  assign n18149 = n18148 ^ n18141;
  assign n18150 = ~n17854 & n18149;
  assign n18151 = n18150 ^ n18148;
  assign n18152 = n17985 ^ n17860;
  assign n18153 = ~n18143 & n18152;
  assign n18154 = n17992 & n18153;
  assign n18155 = ~n18151 & ~n18154;
  assign n18125 = n4040 & ~n10570;
  assign n18126 = x124 & n4267;
  assign n18127 = x126 & n4270;
  assign n18128 = ~n18126 & ~n18127;
  assign n18129 = x125 & n4044;
  assign n18130 = n18128 & ~n18129;
  assign n18131 = ~n18125 & n18130;
  assign n18132 = n18131 ^ x38;
  assign n18115 = n4643 & n9691;
  assign n18116 = x121 & n4653;
  assign n18117 = x123 & n5046;
  assign n18118 = ~n18116 & ~n18117;
  assign n18119 = x122 & n4646;
  assign n18120 = n18118 & ~n18119;
  assign n18121 = ~n18115 & n18120;
  assign n18122 = n18121 ^ x41;
  assign n18103 = n5942 & n7987;
  assign n18104 = x115 & n6186;
  assign n18105 = x117 & n6406;
  assign n18106 = ~n18104 & ~n18105;
  assign n18107 = x116 & n5947;
  assign n18108 = n18106 & ~n18107;
  assign n18109 = ~n18103 & n18108;
  assign n18110 = n18109 ^ x47;
  assign n18092 = n6626 & n7220;
  assign n18093 = x112 & n6884;
  assign n18094 = x113 & n6630;
  assign n18095 = ~n18093 & ~n18094;
  assign n18096 = x114 & n6888;
  assign n18097 = n18095 & ~n18096;
  assign n18098 = ~n18092 & n18097;
  assign n18099 = n18098 ^ x50;
  assign n18089 = n17938 ^ n17927;
  assign n18090 = n17939 & n18089;
  assign n18091 = n18090 ^ n17930;
  assign n18100 = n18099 ^ n18091;
  assign n18079 = n6478 & n7395;
  assign n18080 = x110 & n7400;
  assign n18081 = x109 & n7650;
  assign n18082 = ~n18080 & ~n18081;
  assign n18083 = x111 & n7652;
  assign n18084 = n18082 & ~n18083;
  assign n18085 = ~n18079 & n18084;
  assign n18086 = n18085 ^ x53;
  assign n18076 = n17917 ^ n17914;
  assign n18077 = n17926 & n18076;
  assign n18078 = n18077 ^ n17925;
  assign n18087 = n18086 ^ n18078;
  assign n18066 = n5792 & n8171;
  assign n18067 = x106 & n8181;
  assign n18068 = x107 & n8174;
  assign n18069 = ~n18067 & ~n18068;
  assign n18070 = x108 & n8732;
  assign n18071 = n18069 & ~n18070;
  assign n18072 = ~n18066 & n18071;
  assign n18073 = n18072 ^ x56;
  assign n18063 = n17904 ^ n17883;
  assign n18064 = n17913 & n18063;
  assign n18065 = n18064 ^ n17912;
  assign n18074 = n18073 ^ n18065;
  assign n18054 = n5117 & n9002;
  assign n18055 = x103 & n9012;
  assign n18056 = x104 & n9005;
  assign n18057 = ~n18055 & ~n18056;
  assign n18058 = x105 & n9557;
  assign n18059 = n18057 & ~n18058;
  assign n18060 = ~n18054 & n18059;
  assign n18061 = n18060 ^ x59;
  assign n18049 = n17894 ^ n17886;
  assign n18050 = ~n17903 & ~n18049;
  assign n18051 = n18050 ^ n17902;
  assign n18041 = n3568 ^ x63;
  assign n18042 = n18041 ^ n3568;
  assign n18043 = n3568 ^ n3392;
  assign n18044 = n18043 ^ n3568;
  assign n18045 = n18042 & n18044;
  assign n18046 = n18045 ^ n3568;
  assign n18047 = ~n10177 & n18046;
  assign n18048 = n18047 ^ n3568;
  assign n18052 = n18051 ^ n18048;
  assign n18033 = n4509 & n9878;
  assign n18034 = x100 & n9888;
  assign n18035 = x102 & n10501;
  assign n18036 = ~n18034 & ~n18035;
  assign n18037 = x101 & n9881;
  assign n18038 = n18036 & ~n18037;
  assign n18039 = ~n18033 & n18038;
  assign n18040 = n18039 ^ x62;
  assign n18053 = n18052 ^ n18040;
  assign n18062 = n18061 ^ n18053;
  assign n18075 = n18074 ^ n18062;
  assign n18088 = n18087 ^ n18075;
  assign n18101 = n18100 ^ n18088;
  assign n18030 = n17943 ^ n17940;
  assign n18031 = n17952 & n18030;
  assign n18032 = n18031 ^ n17951;
  assign n18102 = n18101 ^ n18032;
  assign n18111 = n18110 ^ n18102;
  assign n18027 = n17961 ^ n17880;
  assign n18028 = n17962 & n18027;
  assign n18029 = n18028 ^ n17880;
  assign n18112 = n18111 ^ n18029;
  assign n18019 = n5262 & n8820;
  assign n18020 = x118 & n5488;
  assign n18021 = x120 & n5491;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = x119 & n5266;
  assign n18024 = n18022 & ~n18023;
  assign n18025 = ~n18019 & n18024;
  assign n18026 = n18025 ^ x44;
  assign n18113 = n18112 ^ n18026;
  assign n18016 = n17963 ^ n17874;
  assign n18017 = ~n17964 & n18016;
  assign n18018 = n18017 ^ n17877;
  assign n18114 = n18113 ^ n18018;
  assign n18123 = n18122 ^ n18114;
  assign n18013 = n17974 ^ n17866;
  assign n18014 = n17966 & n18013;
  assign n18015 = n18014 ^ n17974;
  assign n18124 = n18123 ^ n18015;
  assign n18133 = n18132 ^ n18124;
  assign n18010 = n17984 ^ n17975;
  assign n18011 = n17976 & ~n18010;
  assign n18012 = n18011 ^ n17984;
  assign n18134 = n18133 ^ n18012;
  assign n17996 = x127 & n3356;
  assign n17997 = ~x35 & ~n17996;
  assign n17998 = n17997 ^ x34;
  assign n17999 = n3175 & n11409;
  assign n18000 = n17999 ^ n17997;
  assign n18001 = ~n17997 & n18000;
  assign n18002 = n18001 ^ n17997;
  assign n18003 = x127 & n3698;
  assign n18004 = ~n18002 & ~n18003;
  assign n18005 = n18004 ^ n18001;
  assign n18006 = n18005 ^ n17997;
  assign n18007 = n18006 ^ n17999;
  assign n18008 = ~n17998 & n18007;
  assign n18009 = n18008 ^ x34;
  assign n18135 = n18134 ^ n18009;
  assign n18156 = n18155 ^ n18135;
  assign n18305 = ~n18135 & ~n18136;
  assign n18306 = ~n18142 & ~n18305;
  assign n18307 = ~n18135 & ~n18144;
  assign n18308 = ~n18137 & ~n18307;
  assign n18309 = ~n18306 & ~n18308;
  assign n18310 = n17854 & ~n18309;
  assign n18311 = n18135 & n18140;
  assign n18312 = n18136 & n18308;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = ~n18310 & n18313;
  assign n18294 = n4040 & ~n10855;
  assign n18295 = x125 & n4267;
  assign n18296 = x127 & n4270;
  assign n18297 = ~n18295 & ~n18296;
  assign n18298 = x126 & n4044;
  assign n18299 = n18297 & ~n18298;
  assign n18300 = ~n18294 & n18299;
  assign n18301 = n18300 ^ x38;
  assign n18284 = n4643 & n9999;
  assign n18285 = x122 & n4653;
  assign n18286 = x123 & n4646;
  assign n18287 = ~n18285 & ~n18286;
  assign n18288 = x124 & n5046;
  assign n18289 = n18287 & ~n18288;
  assign n18290 = ~n18284 & n18289;
  assign n18291 = n18290 ^ x41;
  assign n18274 = n5262 & n9094;
  assign n18275 = x119 & n5488;
  assign n18276 = x121 & n5491;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = x120 & n5266;
  assign n18279 = n18277 & ~n18278;
  assign n18280 = ~n18274 & n18279;
  assign n18281 = n18280 ^ x44;
  assign n18260 = n6728 & n7395;
  assign n18261 = x111 & n7400;
  assign n18262 = x110 & n7650;
  assign n18263 = ~n18261 & ~n18262;
  assign n18264 = x112 & n7652;
  assign n18265 = n18263 & ~n18264;
  assign n18266 = ~n18260 & n18265;
  assign n18267 = n18266 ^ x53;
  assign n18250 = n6026 & n8171;
  assign n18251 = x107 & n8181;
  assign n18252 = x109 & n8732;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = x108 & n8174;
  assign n18255 = n18253 & ~n18254;
  assign n18256 = ~n18250 & n18255;
  assign n18257 = n18256 ^ x56;
  assign n18247 = n18073 ^ n18062;
  assign n18248 = n18074 & n18247;
  assign n18249 = n18248 ^ n18065;
  assign n18258 = n18257 ^ n18249;
  assign n18237 = n5351 & n9002;
  assign n18238 = x104 & n9012;
  assign n18239 = x106 & n9557;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = x105 & n9005;
  assign n18242 = n18240 & ~n18241;
  assign n18243 = ~n18237 & n18242;
  assign n18244 = n18243 ^ x59;
  assign n18234 = n18061 ^ n18052;
  assign n18235 = n18053 & ~n18234;
  assign n18236 = n18235 ^ n18061;
  assign n18245 = n18244 ^ n18236;
  assign n18212 = n17885 ^ x99;
  assign n18213 = n18212 ^ n17885;
  assign n18214 = n17885 ^ n10177;
  assign n18215 = n18214 ^ n17885;
  assign n18216 = ~n18213 & n18215;
  assign n18217 = n18216 ^ n17885;
  assign n18218 = x98 & n18217;
  assign n18219 = n18218 ^ n17885;
  assign n18220 = n18051 & ~n18219;
  assign n18221 = n10177 ^ x98;
  assign n18222 = n3568 ^ x99;
  assign n18223 = n18222 ^ n18221;
  assign n18224 = x97 ^ x63;
  assign n18225 = ~x97 & ~n18224;
  assign n18226 = n18225 ^ x99;
  assign n18227 = n18226 ^ x97;
  assign n18228 = n18223 & ~n18227;
  assign n18229 = n18228 ^ n18225;
  assign n18230 = n18229 ^ x97;
  assign n18231 = n18221 & ~n18230;
  assign n18232 = ~n18220 & ~n18231;
  assign n18203 = n4718 & n9878;
  assign n18204 = x101 & n9888;
  assign n18205 = x103 & n10501;
  assign n18206 = ~n18204 & ~n18205;
  assign n18207 = x102 & n9881;
  assign n18208 = n18206 & ~n18207;
  assign n18209 = ~n18203 & n18208;
  assign n18210 = n18209 ^ x62;
  assign n18194 = n3749 ^ x63;
  assign n18195 = n18194 ^ n3749;
  assign n18196 = n3749 ^ n3568;
  assign n18197 = n18196 ^ n3749;
  assign n18198 = n18195 & n18197;
  assign n18199 = n18198 ^ n3749;
  assign n18200 = ~n10177 & n18199;
  assign n18201 = n18200 ^ n3749;
  assign n18202 = n18201 ^ x35;
  assign n18211 = n18210 ^ n18202;
  assign n18233 = n18232 ^ n18211;
  assign n18246 = n18245 ^ n18233;
  assign n18259 = n18258 ^ n18246;
  assign n18268 = n18267 ^ n18259;
  assign n18191 = n18078 ^ n18075;
  assign n18192 = n18087 & n18191;
  assign n18193 = n18192 ^ n18086;
  assign n18269 = n18268 ^ n18193;
  assign n18188 = n18091 ^ n18088;
  assign n18189 = n18100 & n18188;
  assign n18190 = n18189 ^ n18099;
  assign n18270 = n18269 ^ n18190;
  assign n18180 = n6626 & n7481;
  assign n18181 = x113 & n6884;
  assign n18182 = x115 & n6888;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = x114 & n6630;
  assign n18185 = n18183 & ~n18184;
  assign n18186 = ~n18180 & n18185;
  assign n18187 = n18186 ^ x50;
  assign n18271 = n18270 ^ n18187;
  assign n18172 = n5942 & n8265;
  assign n18173 = x116 & n6186;
  assign n18174 = x117 & n5947;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = x118 & n6406;
  assign n18177 = n18175 & ~n18176;
  assign n18178 = ~n18172 & n18177;
  assign n18179 = n18178 ^ x47;
  assign n18272 = n18271 ^ n18179;
  assign n18169 = n18110 ^ n18101;
  assign n18170 = n18102 & ~n18169;
  assign n18171 = n18170 ^ n18110;
  assign n18273 = n18272 ^ n18171;
  assign n18282 = n18281 ^ n18273;
  assign n18166 = n18111 ^ n18026;
  assign n18167 = ~n18112 & n18166;
  assign n18168 = n18167 ^ n18029;
  assign n18283 = n18282 ^ n18168;
  assign n18292 = n18291 ^ n18283;
  assign n18163 = n18122 ^ n18018;
  assign n18164 = n18114 & n18163;
  assign n18165 = n18164 ^ n18122;
  assign n18293 = n18292 ^ n18165;
  assign n18302 = n18301 ^ n18293;
  assign n18160 = n18132 ^ n18123;
  assign n18161 = n18124 & ~n18160;
  assign n18162 = n18161 ^ n18132;
  assign n18303 = n18302 ^ n18162;
  assign n18157 = n18133 ^ n18009;
  assign n18158 = n18134 & n18157;
  assign n18159 = n18158 ^ n18009;
  assign n18304 = n18303 ^ n18159;
  assign n18315 = n18314 ^ n18304;
  assign n18433 = n4643 & n10303;
  assign n18434 = x123 & n4653;
  assign n18435 = x124 & n4646;
  assign n18436 = ~n18434 & ~n18435;
  assign n18437 = x125 & n5046;
  assign n18438 = n18436 & ~n18437;
  assign n18439 = ~n18433 & n18438;
  assign n18440 = n18439 ^ x41;
  assign n18423 = n5262 & n9387;
  assign n18424 = x120 & n5488;
  assign n18425 = x121 & n5266;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = x122 & n5491;
  assign n18428 = n18426 & ~n18427;
  assign n18429 = ~n18423 & n18428;
  assign n18430 = n18429 ^ x44;
  assign n18410 = n6626 & n7730;
  assign n18411 = x114 & n6884;
  assign n18412 = x116 & n6888;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = x115 & n6630;
  assign n18415 = n18413 & ~n18414;
  assign n18416 = ~n18410 & n18415;
  assign n18417 = n18416 ^ x50;
  assign n18407 = n18267 ^ n18193;
  assign n18408 = n18268 & n18407;
  assign n18409 = n18408 ^ n18193;
  assign n18418 = n18417 ^ n18409;
  assign n18397 = n6975 & n7395;
  assign n18398 = x111 & n7650;
  assign n18399 = x112 & n7400;
  assign n18400 = ~n18398 & ~n18399;
  assign n18401 = x113 & n7652;
  assign n18402 = n18400 & ~n18401;
  assign n18403 = ~n18397 & n18402;
  assign n18404 = n18403 ^ x53;
  assign n18394 = n18257 ^ n18246;
  assign n18395 = n18258 & n18394;
  assign n18396 = n18395 ^ n18249;
  assign n18405 = n18404 ^ n18396;
  assign n18384 = n6250 & n8171;
  assign n18385 = x108 & n8181;
  assign n18386 = x110 & n8732;
  assign n18387 = ~n18385 & ~n18386;
  assign n18388 = x109 & n8174;
  assign n18389 = n18387 & ~n18388;
  assign n18390 = ~n18384 & n18389;
  assign n18391 = n18390 ^ x56;
  assign n18381 = n18244 ^ n18233;
  assign n18382 = n18245 & n18381;
  assign n18383 = n18382 ^ n18236;
  assign n18392 = n18391 ^ n18383;
  assign n18371 = n5578 & n9002;
  assign n18372 = x105 & n9012;
  assign n18373 = x106 & n9005;
  assign n18374 = ~n18372 & ~n18373;
  assign n18375 = x107 & n9557;
  assign n18376 = n18374 & ~n18375;
  assign n18377 = ~n18371 & n18376;
  assign n18378 = n18377 ^ x59;
  assign n18368 = n18232 ^ n18210;
  assign n18369 = ~n18211 & ~n18368;
  assign n18370 = n18369 ^ n18232;
  assign n18379 = n18378 ^ n18370;
  assign n18359 = n4912 & n9878;
  assign n18360 = x102 & n9888;
  assign n18361 = x103 & n9881;
  assign n18362 = ~n18360 & ~n18361;
  assign n18363 = x104 & n10501;
  assign n18364 = n18362 & ~n18363;
  assign n18365 = ~n18359 & n18364;
  assign n18366 = n18365 ^ x62;
  assign n18355 = x101 & n10177;
  assign n18356 = x100 & n12123;
  assign n18357 = ~n18355 & ~n18356;
  assign n18348 = x99 ^ x35;
  assign n18349 = n3750 & ~n12123;
  assign n18350 = n18349 ^ x98;
  assign n18351 = n18350 ^ x99;
  assign n18352 = ~n18348 & n18351;
  assign n18353 = n18352 ^ x99;
  assign n18354 = ~n12893 & n18353;
  assign n18358 = n18357 ^ n18354;
  assign n18367 = n18366 ^ n18358;
  assign n18380 = n18379 ^ n18367;
  assign n18393 = n18392 ^ n18380;
  assign n18406 = n18405 ^ n18393;
  assign n18419 = n18418 ^ n18406;
  assign n18345 = n18269 ^ n18187;
  assign n18346 = ~n18270 & n18345;
  assign n18347 = n18346 ^ n18190;
  assign n18420 = n18419 ^ n18347;
  assign n18337 = n5942 & n8542;
  assign n18338 = x117 & n6186;
  assign n18339 = x118 & n5947;
  assign n18340 = ~n18338 & ~n18339;
  assign n18341 = x119 & n6406;
  assign n18342 = n18340 & ~n18341;
  assign n18343 = ~n18337 & n18342;
  assign n18344 = n18343 ^ x47;
  assign n18421 = n18420 ^ n18344;
  assign n18334 = n18179 ^ n18171;
  assign n18335 = ~n18272 & ~n18334;
  assign n18336 = n18335 ^ n18271;
  assign n18422 = n18421 ^ n18336;
  assign n18431 = n18430 ^ n18422;
  assign n18331 = n18281 ^ n18168;
  assign n18332 = n18282 & n18331;
  assign n18333 = n18332 ^ n18168;
  assign n18432 = n18431 ^ n18333;
  assign n18441 = n18440 ^ n18432;
  assign n18328 = n18291 ^ n18165;
  assign n18329 = n18292 & n18328;
  assign n18330 = n18329 ^ n18165;
  assign n18442 = n18441 ^ n18330;
  assign n18322 = n4040 & ~n10281;
  assign n18323 = x126 & n4267;
  assign n18324 = x127 & n4044;
  assign n18325 = ~n18323 & ~n18324;
  assign n18326 = ~n18322 & n18325;
  assign n18327 = n18326 ^ x38;
  assign n18443 = n18442 ^ n18327;
  assign n18319 = n18301 ^ n18162;
  assign n18320 = n18302 & n18319;
  assign n18321 = n18320 ^ n18162;
  assign n18444 = n18443 ^ n18321;
  assign n18316 = n18314 ^ n18159;
  assign n18317 = ~n18304 & n18316;
  assign n18318 = n18317 ^ n18314;
  assign n18445 = n18444 ^ n18318;
  assign n18579 = n4643 & ~n10570;
  assign n18580 = x124 & n4653;
  assign n18581 = x125 & n4646;
  assign n18582 = ~n18580 & ~n18581;
  assign n18583 = x126 & n5046;
  assign n18584 = n18582 & ~n18583;
  assign n18585 = ~n18579 & n18584;
  assign n18586 = n18585 ^ x41;
  assign n18569 = n5262 & n9691;
  assign n18570 = x121 & n5488;
  assign n18571 = x122 & n5266;
  assign n18572 = ~n18570 & ~n18571;
  assign n18573 = x123 & n5491;
  assign n18574 = n18572 & ~n18573;
  assign n18575 = ~n18569 & n18574;
  assign n18576 = n18575 ^ x44;
  assign n18556 = n6626 & n7987;
  assign n18557 = x115 & n6884;
  assign n18558 = x117 & n6888;
  assign n18559 = ~n18557 & ~n18558;
  assign n18560 = x116 & n6630;
  assign n18561 = n18559 & ~n18560;
  assign n18562 = ~n18556 & n18561;
  assign n18563 = n18562 ^ x50;
  assign n18547 = n7220 & n7395;
  assign n18548 = x112 & n7650;
  assign n18549 = x113 & n7400;
  assign n18550 = ~n18548 & ~n18549;
  assign n18551 = x114 & n7652;
  assign n18552 = n18550 & ~n18551;
  assign n18553 = ~n18547 & n18552;
  assign n18554 = n18553 ^ x53;
  assign n18536 = n6478 & n8171;
  assign n18537 = x109 & n8181;
  assign n18538 = x110 & n8174;
  assign n18539 = ~n18537 & ~n18538;
  assign n18540 = x111 & n8732;
  assign n18541 = n18539 & ~n18540;
  assign n18542 = ~n18536 & n18541;
  assign n18543 = n18542 ^ x56;
  assign n18533 = n18378 ^ n18367;
  assign n18534 = ~n18379 & ~n18533;
  assign n18535 = n18534 ^ n18370;
  assign n18544 = n18543 ^ n18535;
  assign n18523 = n5792 & n9002;
  assign n18524 = x107 & n9005;
  assign n18525 = x106 & n9012;
  assign n18526 = ~n18524 & ~n18525;
  assign n18527 = x108 & n9557;
  assign n18528 = n18526 & ~n18527;
  assign n18529 = ~n18523 & n18528;
  assign n18530 = n18529 ^ x59;
  assign n18503 = n18356 ^ x102;
  assign n18504 = n18503 ^ n18356;
  assign n18505 = n18356 ^ n10177;
  assign n18506 = n18505 ^ n18356;
  assign n18507 = ~n18504 & n18506;
  assign n18508 = n18507 ^ n18356;
  assign n18509 = x101 & n18508;
  assign n18510 = n18509 ^ n18356;
  assign n18512 = ~x101 & x102;
  assign n18511 = ~x100 & x101;
  assign n18513 = n18512 ^ n18511;
  assign n18514 = n18513 ^ n18512;
  assign n18515 = n18512 ^ x63;
  assign n18516 = n18515 ^ n18512;
  assign n18517 = n18514 & n18516;
  assign n18518 = n18517 ^ n18512;
  assign n18519 = ~n10177 & n18518;
  assign n18520 = n18519 ^ n18512;
  assign n18521 = ~n18510 & ~n18520;
  assign n18500 = n18366 ^ n18354;
  assign n18501 = ~n18358 & ~n18500;
  assign n18502 = n18501 ^ n18366;
  assign n18522 = n18521 ^ n18502;
  assign n18531 = n18530 ^ n18522;
  assign n18492 = n5117 & n9878;
  assign n18493 = x104 & n9881;
  assign n18494 = x103 & n9888;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = x105 & n10501;
  assign n18497 = n18495 & ~n18496;
  assign n18498 = ~n18492 & n18497;
  assign n18499 = n18498 ^ x62;
  assign n18532 = n18531 ^ n18499;
  assign n18545 = n18544 ^ n18532;
  assign n18489 = n18391 ^ n18380;
  assign n18490 = n18392 & n18489;
  assign n18491 = n18490 ^ n18383;
  assign n18546 = n18545 ^ n18491;
  assign n18555 = n18554 ^ n18546;
  assign n18564 = n18563 ^ n18555;
  assign n18486 = n18396 ^ n18393;
  assign n18487 = n18405 & n18486;
  assign n18488 = n18487 ^ n18404;
  assign n18565 = n18564 ^ n18488;
  assign n18483 = n18409 ^ n18406;
  assign n18484 = n18418 & n18483;
  assign n18485 = n18484 ^ n18417;
  assign n18566 = n18565 ^ n18485;
  assign n18475 = n5942 & n8820;
  assign n18476 = x118 & n6186;
  assign n18477 = x119 & n5947;
  assign n18478 = ~n18476 & ~n18477;
  assign n18479 = x120 & n6406;
  assign n18480 = n18478 & ~n18479;
  assign n18481 = ~n18475 & n18480;
  assign n18482 = n18481 ^ x47;
  assign n18567 = n18566 ^ n18482;
  assign n18472 = n18419 ^ n18344;
  assign n18473 = ~n18420 & n18472;
  assign n18474 = n18473 ^ n18347;
  assign n18568 = n18567 ^ n18474;
  assign n18577 = n18576 ^ n18568;
  assign n18469 = n18430 ^ n18336;
  assign n18470 = ~n18422 & ~n18469;
  assign n18471 = n18470 ^ n18430;
  assign n18578 = n18577 ^ n18471;
  assign n18587 = n18586 ^ n18578;
  assign n18466 = n18440 ^ n18333;
  assign n18467 = ~n18432 & n18466;
  assign n18468 = n18467 ^ n18440;
  assign n18588 = n18587 ^ n18468;
  assign n18452 = x127 & n3879;
  assign n18453 = ~x38 & ~n18452;
  assign n18454 = n18453 ^ x37;
  assign n18455 = n3693 & n11409;
  assign n18456 = n18455 ^ n18453;
  assign n18457 = ~n18453 & n18456;
  assign n18458 = n18457 ^ n18453;
  assign n18459 = x127 & n4266;
  assign n18460 = ~n18458 & ~n18459;
  assign n18461 = n18460 ^ n18457;
  assign n18462 = n18461 ^ n18453;
  assign n18463 = n18462 ^ n18455;
  assign n18464 = ~n18454 & n18463;
  assign n18465 = n18464 ^ x37;
  assign n18589 = n18588 ^ n18465;
  assign n18449 = n18441 ^ n18327;
  assign n18450 = n18442 & ~n18449;
  assign n18451 = n18450 ^ n18330;
  assign n18590 = n18589 ^ n18451;
  assign n18446 = n18321 ^ n18318;
  assign n18447 = ~n18444 & ~n18446;
  assign n18448 = n18447 ^ n18318;
  assign n18591 = n18590 ^ n18448;
  assign n18709 = n18451 ^ n18448;
  assign n18710 = ~n18590 & ~n18709;
  assign n18711 = n18710 ^ n18448;
  assign n18693 = n6626 & n8265;
  assign n18694 = x116 & n6884;
  assign n18695 = x118 & n6888;
  assign n18696 = ~n18694 & ~n18695;
  assign n18697 = x117 & n6630;
  assign n18698 = n18696 & ~n18697;
  assign n18699 = ~n18693 & n18698;
  assign n18700 = n18699 ^ x50;
  assign n18690 = n18555 ^ n18488;
  assign n18691 = ~n18564 & n18690;
  assign n18692 = n18691 ^ n18563;
  assign n18701 = n18700 ^ n18692;
  assign n18680 = n7395 & n7481;
  assign n18681 = x113 & n7650;
  assign n18682 = x114 & n7400;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = x115 & n7652;
  assign n18685 = n18683 & ~n18684;
  assign n18686 = ~n18680 & n18685;
  assign n18687 = n18686 ^ x53;
  assign n18677 = n18554 ^ n18491;
  assign n18678 = n18546 & n18677;
  assign n18679 = n18678 ^ n18554;
  assign n18688 = n18687 ^ n18679;
  assign n18667 = n6728 & n8171;
  assign n18668 = x110 & n8181;
  assign n18669 = x111 & n8174;
  assign n18670 = ~n18668 & ~n18669;
  assign n18671 = x112 & n8732;
  assign n18672 = n18670 & ~n18671;
  assign n18673 = ~n18667 & n18672;
  assign n18674 = n18673 ^ x56;
  assign n18664 = n18535 ^ n18532;
  assign n18665 = ~n18544 & n18664;
  assign n18666 = n18665 ^ n18543;
  assign n18675 = n18674 ^ n18666;
  assign n18654 = n6026 & n9002;
  assign n18655 = x107 & n9012;
  assign n18656 = x109 & n9557;
  assign n18657 = ~n18655 & ~n18656;
  assign n18658 = x108 & n9005;
  assign n18659 = n18657 & ~n18658;
  assign n18660 = ~n18654 & n18659;
  assign n18661 = n18660 ^ x59;
  assign n18651 = n18522 ^ n18499;
  assign n18652 = n18531 & ~n18651;
  assign n18653 = n18652 ^ n18530;
  assign n18662 = n18661 ^ n18653;
  assign n18641 = n5351 & n9878;
  assign n18642 = x104 & n9888;
  assign n18643 = x106 & n10501;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = x105 & n9881;
  assign n18646 = n18644 & ~n18645;
  assign n18647 = ~n18641 & n18646;
  assign n18648 = n18647 ^ x62;
  assign n18631 = x103 ^ x102;
  assign n18632 = n18631 ^ x103;
  assign n18633 = x103 ^ x63;
  assign n18634 = n18633 ^ x103;
  assign n18635 = n18632 & n18634;
  assign n18636 = n18635 ^ x103;
  assign n18637 = ~n10177 & n18636;
  assign n18638 = n18637 ^ x103;
  assign n18639 = n18638 ^ n18357;
  assign n18640 = n18639 ^ x38;
  assign n18649 = n18648 ^ n18640;
  assign n18629 = n18502 & n18521;
  assign n18630 = n18629 ^ n18510;
  assign n18650 = n18649 ^ n18630;
  assign n18663 = n18662 ^ n18650;
  assign n18676 = n18675 ^ n18663;
  assign n18689 = n18688 ^ n18676;
  assign n18702 = n18701 ^ n18689;
  assign n18621 = n5942 & n9094;
  assign n18622 = x119 & n6186;
  assign n18623 = x120 & n5947;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 = x121 & n6406;
  assign n18626 = n18624 & ~n18625;
  assign n18627 = ~n18621 & n18626;
  assign n18628 = n18627 ^ x47;
  assign n18703 = n18702 ^ n18628;
  assign n18618 = n18485 ^ n18482;
  assign n18619 = ~n18566 & ~n18618;
  assign n18620 = n18619 ^ n18565;
  assign n18704 = n18703 ^ n18620;
  assign n18615 = n18576 ^ n18474;
  assign n18616 = n18568 & n18615;
  assign n18617 = n18616 ^ n18576;
  assign n18705 = n18704 ^ n18617;
  assign n18607 = n5262 & n9999;
  assign n18608 = x122 & n5488;
  assign n18609 = x123 & n5266;
  assign n18610 = ~n18608 & ~n18609;
  assign n18611 = x124 & n5491;
  assign n18612 = n18610 & ~n18611;
  assign n18613 = ~n18607 & n18612;
  assign n18614 = n18613 ^ x44;
  assign n18706 = n18705 ^ n18614;
  assign n18604 = n18587 ^ n18465;
  assign n18605 = n18588 & n18604;
  assign n18606 = n18605 ^ n18465;
  assign n18707 = n18706 ^ n18606;
  assign n18595 = n4643 & ~n10855;
  assign n18596 = x125 & n4653;
  assign n18597 = x127 & n5046;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = x126 & n4646;
  assign n18600 = n18598 & ~n18599;
  assign n18601 = ~n18595 & n18600;
  assign n18602 = n18601 ^ x41;
  assign n18592 = n18586 ^ n18471;
  assign n18593 = n18578 & n18592;
  assign n18594 = n18593 ^ n18586;
  assign n18603 = n18602 ^ n18594;
  assign n18708 = n18707 ^ n18603;
  assign n18712 = n18711 ^ n18708;
  assign n18824 = n18594 & n18602;
  assign n18823 = ~n18594 & ~n18602;
  assign n18825 = n18824 ^ n18823;
  assign n18826 = ~n18706 & n18825;
  assign n18827 = n18826 ^ n18824;
  assign n18828 = n18707 & n18827;
  assign n18842 = n18824 ^ n18706;
  assign n18843 = ~n18707 & ~n18842;
  assign n18844 = n18843 ^ n18606;
  assign n18845 = ~n18823 & ~n18844;
  assign n18829 = n18706 ^ n18603;
  assign n18830 = n18829 ^ n18707;
  assign n18831 = n18606 ^ n18602;
  assign n18832 = n18831 ^ n18706;
  assign n18833 = n18832 ^ n18706;
  assign n18834 = ~n18603 & ~n18833;
  assign n18835 = n18834 ^ n18603;
  assign n18836 = ~n18832 & ~n18835;
  assign n18837 = n18836 ^ n18706;
  assign n18838 = ~n18830 & n18837;
  assign n18839 = n18838 ^ n18834;
  assign n18840 = n18839 ^ n18706;
  assign n18841 = n18840 ^ n18707;
  assign n18846 = n18845 ^ n18841;
  assign n18847 = ~n18711 & n18846;
  assign n18848 = n18847 ^ n18841;
  assign n18849 = ~n18828 & ~n18848;
  assign n18811 = n5262 & n10303;
  assign n18812 = x123 & n5488;
  assign n18813 = x124 & n5266;
  assign n18814 = ~n18812 & ~n18813;
  assign n18815 = x125 & n5491;
  assign n18816 = n18814 & ~n18815;
  assign n18817 = ~n18811 & n18816;
  assign n18818 = n18817 ^ x44;
  assign n18801 = n5942 & n9387;
  assign n18802 = x120 & n6186;
  assign n18803 = x122 & n6406;
  assign n18804 = ~n18802 & ~n18803;
  assign n18805 = x121 & n5947;
  assign n18806 = n18804 & ~n18805;
  assign n18807 = ~n18801 & n18806;
  assign n18808 = n18807 ^ x47;
  assign n18791 = n6626 & n8542;
  assign n18792 = x117 & n6884;
  assign n18793 = x118 & n6630;
  assign n18794 = ~n18792 & ~n18793;
  assign n18795 = x119 & n6888;
  assign n18796 = n18794 & ~n18795;
  assign n18797 = ~n18791 & n18796;
  assign n18798 = n18797 ^ x50;
  assign n18781 = n7395 & n7730;
  assign n18782 = x114 & n7650;
  assign n18783 = x115 & n7400;
  assign n18784 = ~n18782 & ~n18783;
  assign n18785 = x116 & n7652;
  assign n18786 = n18784 & ~n18785;
  assign n18787 = ~n18781 & n18786;
  assign n18788 = n18787 ^ x53;
  assign n18778 = n18674 ^ n18663;
  assign n18779 = n18675 & n18778;
  assign n18780 = n18779 ^ n18666;
  assign n18789 = n18788 ^ n18780;
  assign n18768 = n6975 & n8171;
  assign n18769 = x111 & n8181;
  assign n18770 = x113 & n8732;
  assign n18771 = ~n18769 & ~n18770;
  assign n18772 = x112 & n8174;
  assign n18773 = n18771 & ~n18772;
  assign n18774 = ~n18768 & n18773;
  assign n18775 = n18774 ^ x56;
  assign n18765 = n18661 ^ n18650;
  assign n18766 = n18662 & n18765;
  assign n18767 = n18766 ^ n18653;
  assign n18776 = n18775 ^ n18767;
  assign n18755 = n6250 & n9002;
  assign n18756 = x108 & n9012;
  assign n18757 = x109 & n9005;
  assign n18758 = ~n18756 & ~n18757;
  assign n18759 = x110 & n9557;
  assign n18760 = n18758 & ~n18759;
  assign n18761 = ~n18755 & n18760;
  assign n18762 = n18761 ^ x59;
  assign n18746 = n5578 & n9878;
  assign n18747 = x105 & n9888;
  assign n18748 = x107 & n10501;
  assign n18749 = ~n18747 & ~n18748;
  assign n18750 = x106 & n9881;
  assign n18751 = n18749 & ~n18750;
  assign n18752 = ~n18746 & n18751;
  assign n18753 = n18752 ^ x62;
  assign n18742 = n18357 ^ x38;
  assign n18743 = n18639 & n18742;
  assign n18744 = n18743 ^ x38;
  assign n18734 = x104 ^ x63;
  assign n18735 = n18734 ^ x104;
  assign n18736 = x104 ^ x103;
  assign n18737 = n18736 ^ x104;
  assign n18738 = n18735 & n18737;
  assign n18739 = n18738 ^ x104;
  assign n18740 = ~n10177 & n18739;
  assign n18741 = n18740 ^ x104;
  assign n18745 = n18744 ^ n18741;
  assign n18754 = n18753 ^ n18745;
  assign n18763 = n18762 ^ n18754;
  assign n18731 = n18648 ^ n18630;
  assign n18732 = n18649 & n18731;
  assign n18733 = n18732 ^ n18630;
  assign n18764 = n18763 ^ n18733;
  assign n18777 = n18776 ^ n18764;
  assign n18790 = n18789 ^ n18777;
  assign n18799 = n18798 ^ n18790;
  assign n18728 = n18687 ^ n18676;
  assign n18729 = n18688 & n18728;
  assign n18730 = n18729 ^ n18679;
  assign n18800 = n18799 ^ n18730;
  assign n18809 = n18808 ^ n18800;
  assign n18725 = n18700 ^ n18689;
  assign n18726 = n18701 & n18725;
  assign n18727 = n18726 ^ n18692;
  assign n18810 = n18809 ^ n18727;
  assign n18819 = n18818 ^ n18810;
  assign n18722 = n18628 ^ n18620;
  assign n18723 = ~n18703 & n18722;
  assign n18724 = n18723 ^ n18702;
  assign n18820 = n18819 ^ n18724;
  assign n18719 = n18704 ^ n18614;
  assign n18720 = n18705 & ~n18719;
  assign n18721 = n18720 ^ n18617;
  assign n18821 = n18820 ^ n18721;
  assign n18713 = n4643 & ~n10281;
  assign n18714 = x126 & n4653;
  assign n18715 = x127 & n4646;
  assign n18716 = ~n18714 & ~n18715;
  assign n18717 = ~n18713 & n18716;
  assign n18718 = n18717 ^ x41;
  assign n18822 = n18821 ^ n18718;
  assign n18850 = n18849 ^ n18822;
  assign n18958 = n18606 & ~n18706;
  assign n18959 = ~n18822 & ~n18958;
  assign n18960 = n18711 ^ n18602;
  assign n18961 = n18603 & n18960;
  assign n18962 = n18961 ^ n18594;
  assign n18963 = ~n18959 & ~n18962;
  assign n18964 = ~n18606 & n18706;
  assign n18965 = ~n18822 & ~n18823;
  assign n18966 = ~n18964 & ~n18965;
  assign n18967 = n18711 & n18966;
  assign n18968 = n18822 & n18844;
  assign n18969 = ~n18967 & ~n18968;
  assign n18970 = ~n18963 & n18969;
  assign n18951 = n4643 & n11409;
  assign n18952 = x127 & n4653;
  assign n18953 = ~n18951 & ~n18952;
  assign n18954 = n18953 ^ x41;
  assign n18948 = n18810 ^ n18724;
  assign n18949 = n18819 & n18948;
  assign n18950 = n18949 ^ n18818;
  assign n18955 = n18954 ^ n18950;
  assign n18939 = n5262 & ~n10570;
  assign n18940 = x125 & n5266;
  assign n18941 = x124 & n5488;
  assign n18942 = ~n18940 & ~n18941;
  assign n18943 = x126 & n5491;
  assign n18944 = n18942 & ~n18943;
  assign n18945 = ~n18939 & n18944;
  assign n18946 = n18945 ^ x44;
  assign n18926 = n6626 & n8820;
  assign n18927 = x118 & n6884;
  assign n18928 = x119 & n6630;
  assign n18929 = ~n18927 & ~n18928;
  assign n18930 = x120 & n6888;
  assign n18931 = n18929 & ~n18930;
  assign n18932 = ~n18926 & n18931;
  assign n18933 = n18932 ^ x50;
  assign n18923 = n18788 ^ n18777;
  assign n18924 = n18789 & ~n18923;
  assign n18925 = n18924 ^ n18780;
  assign n18934 = n18933 ^ n18925;
  assign n18913 = n7395 & n7987;
  assign n18914 = x115 & n7650;
  assign n18915 = x116 & n7400;
  assign n18916 = ~n18914 & ~n18915;
  assign n18917 = x117 & n7652;
  assign n18918 = n18916 & ~n18917;
  assign n18919 = ~n18913 & n18918;
  assign n18920 = n18919 ^ x53;
  assign n18910 = n18767 ^ n18764;
  assign n18911 = n18776 & ~n18910;
  assign n18912 = n18911 ^ n18775;
  assign n18921 = n18920 ^ n18912;
  assign n18900 = n7220 & n8171;
  assign n18901 = x112 & n8181;
  assign n18902 = x114 & n8732;
  assign n18903 = ~n18901 & ~n18902;
  assign n18904 = x113 & n8174;
  assign n18905 = n18903 & ~n18904;
  assign n18906 = ~n18900 & n18905;
  assign n18907 = n18906 ^ x56;
  assign n18897 = n18762 ^ n18733;
  assign n18898 = ~n18763 & n18897;
  assign n18899 = n18898 ^ n18733;
  assign n18908 = n18907 ^ n18899;
  assign n18888 = n6478 & n9002;
  assign n18889 = x109 & n9012;
  assign n18890 = x110 & n9005;
  assign n18891 = ~n18889 & ~n18890;
  assign n18892 = x111 & n9557;
  assign n18893 = n18891 & ~n18892;
  assign n18894 = ~n18888 & n18893;
  assign n18895 = n18894 ^ x59;
  assign n18878 = x105 ^ x104;
  assign n18879 = n18878 ^ x105;
  assign n18880 = x105 ^ x63;
  assign n18881 = n18880 ^ x105;
  assign n18882 = n18879 & n18881;
  assign n18883 = n18882 ^ x105;
  assign n18884 = ~n10177 & n18883;
  assign n18885 = n18884 ^ x105;
  assign n18876 = n18753 ^ n18744;
  assign n18877 = n18745 & ~n18876;
  assign n18886 = n18885 ^ n18877;
  assign n18868 = n5792 & n9878;
  assign n18869 = x106 & n9888;
  assign n18870 = x108 & n10501;
  assign n18871 = ~n18869 & ~n18870;
  assign n18872 = x107 & n9881;
  assign n18873 = n18871 & ~n18872;
  assign n18874 = ~n18868 & n18873;
  assign n18875 = n18874 ^ x62;
  assign n18887 = n18886 ^ n18875;
  assign n18896 = n18895 ^ n18887;
  assign n18909 = n18908 ^ n18896;
  assign n18922 = n18921 ^ n18909;
  assign n18935 = n18934 ^ n18922;
  assign n18865 = n18790 ^ n18730;
  assign n18866 = n18799 & ~n18865;
  assign n18867 = n18866 ^ n18798;
  assign n18936 = n18935 ^ n18867;
  assign n18857 = n5942 & n9691;
  assign n18858 = x121 & n6186;
  assign n18859 = x123 & n6406;
  assign n18860 = ~n18858 & ~n18859;
  assign n18861 = x122 & n5947;
  assign n18862 = n18860 & ~n18861;
  assign n18863 = ~n18857 & n18862;
  assign n18864 = n18863 ^ x47;
  assign n18937 = n18936 ^ n18864;
  assign n18854 = n18800 ^ n18727;
  assign n18855 = n18809 & ~n18854;
  assign n18856 = n18855 ^ n18808;
  assign n18938 = n18937 ^ n18856;
  assign n18947 = n18946 ^ n18938;
  assign n18956 = n18955 ^ n18947;
  assign n18851 = n18820 ^ n18718;
  assign n18852 = ~n18821 & n18851;
  assign n18853 = n18852 ^ n18721;
  assign n18957 = n18956 ^ n18853;
  assign n18971 = n18970 ^ n18957;
  assign n19083 = n5262 & ~n10855;
  assign n19084 = x125 & n5488;
  assign n19085 = x127 & n5491;
  assign n19086 = ~n19084 & ~n19085;
  assign n19087 = x126 & n5266;
  assign n19088 = n19086 & ~n19087;
  assign n19089 = ~n19083 & n19088;
  assign n19090 = n19089 ^ x44;
  assign n19073 = n5942 & n9999;
  assign n19074 = x122 & n6186;
  assign n19075 = x124 & n6406;
  assign n19076 = ~n19074 & ~n19075;
  assign n19077 = x123 & n5947;
  assign n19078 = n19076 & ~n19077;
  assign n19079 = ~n19073 & n19078;
  assign n19080 = n19079 ^ x47;
  assign n19063 = n6626 & n9094;
  assign n19064 = x120 & n6630;
  assign n19065 = x119 & n6884;
  assign n19066 = ~n19064 & ~n19065;
  assign n19067 = x121 & n6888;
  assign n19068 = n19066 & ~n19067;
  assign n19069 = ~n19063 & n19068;
  assign n19070 = n19069 ^ x50;
  assign n19060 = n18933 ^ n18922;
  assign n19061 = n18934 & n19060;
  assign n19062 = n19061 ^ n18925;
  assign n19071 = n19070 ^ n19062;
  assign n19050 = n7395 & n8265;
  assign n19051 = x116 & n7650;
  assign n19052 = x118 & n7652;
  assign n19053 = ~n19051 & ~n19052;
  assign n19054 = x117 & n7400;
  assign n19055 = n19053 & ~n19054;
  assign n19056 = ~n19050 & n19055;
  assign n19057 = n19056 ^ x53;
  assign n19047 = n18912 ^ n18909;
  assign n19048 = n18921 & n19047;
  assign n19049 = n19048 ^ n18920;
  assign n19058 = n19057 ^ n19049;
  assign n19037 = n7481 & n8171;
  assign n19038 = x113 & n8181;
  assign n19039 = x115 & n8732;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = x114 & n8174;
  assign n19042 = n19040 & ~n19041;
  assign n19043 = ~n19037 & n19042;
  assign n19044 = n19043 ^ x56;
  assign n19027 = n6728 & n9002;
  assign n19028 = x110 & n9012;
  assign n19029 = x111 & n9005;
  assign n19030 = ~n19028 & ~n19029;
  assign n19031 = x112 & n9557;
  assign n19032 = n19030 & ~n19031;
  assign n19033 = ~n19027 & n19032;
  assign n19034 = n19033 ^ x59;
  assign n19017 = n6026 & n9878;
  assign n19018 = x107 & n9888;
  assign n19019 = x109 & n10501;
  assign n19020 = ~n19018 & ~n19019;
  assign n19021 = x108 & n9881;
  assign n19022 = n19020 & ~n19021;
  assign n19023 = ~n19017 & n19022;
  assign n19024 = n19023 ^ x62;
  assign n19014 = n18885 ^ n18741;
  assign n19015 = n18877 & ~n19014;
  assign n19016 = n19015 ^ n18741;
  assign n19025 = n19024 ^ n19016;
  assign n19004 = x106 ^ x63;
  assign n19005 = n19004 ^ x106;
  assign n19006 = x106 ^ x105;
  assign n19007 = n19006 ^ x106;
  assign n19008 = n19005 & n19007;
  assign n19009 = n19008 ^ x106;
  assign n19010 = ~n10177 & n19009;
  assign n19011 = n19010 ^ x106;
  assign n19012 = n19011 ^ n18741;
  assign n19013 = n19012 ^ x41;
  assign n19026 = n19025 ^ n19013;
  assign n19035 = n19034 ^ n19026;
  assign n19001 = n18895 ^ n18886;
  assign n19002 = n18887 & ~n19001;
  assign n19003 = n19002 ^ n18895;
  assign n19036 = n19035 ^ n19003;
  assign n19045 = n19044 ^ n19036;
  assign n18998 = n18899 ^ n18896;
  assign n18999 = n18908 & n18998;
  assign n19000 = n18999 ^ n18907;
  assign n19046 = n19045 ^ n19000;
  assign n19059 = n19058 ^ n19046;
  assign n19072 = n19071 ^ n19059;
  assign n19081 = n19080 ^ n19072;
  assign n18995 = n18935 ^ n18864;
  assign n18996 = ~n18936 & n18995;
  assign n18997 = n18996 ^ n18867;
  assign n19082 = n19081 ^ n18997;
  assign n19091 = n19090 ^ n19082;
  assign n18992 = n18946 ^ n18856;
  assign n18993 = n18938 & n18992;
  assign n18994 = n18993 ^ n18946;
  assign n19092 = n19091 ^ n18994;
  assign n18972 = ~n18947 & n18954;
  assign n18973 = n18950 & n18972;
  assign n18974 = n18853 & n18973;
  assign n18975 = n18947 & ~n18954;
  assign n18976 = ~n18950 & n18975;
  assign n18977 = ~n18853 & n18976;
  assign n18978 = ~n18974 & ~n18977;
  assign n18979 = n18954 ^ n18947;
  assign n18980 = n18955 & n18979;
  assign n18981 = n18980 ^ n18950;
  assign n18982 = n18853 & n18981;
  assign n18983 = ~n18973 & ~n18982;
  assign n18984 = n18983 ^ n18970;
  assign n18985 = n18984 ^ n18983;
  assign n18986 = n18853 & ~n18976;
  assign n18987 = ~n18981 & ~n18986;
  assign n18988 = n18987 ^ n18983;
  assign n18989 = ~n18985 & ~n18988;
  assign n18990 = n18989 ^ n18983;
  assign n18991 = n18978 & n18990;
  assign n19093 = n19092 ^ n18991;
  assign n19194 = ~n18987 & n19092;
  assign n19195 = ~n18974 & ~n19194;
  assign n19196 = ~n18970 & n19195;
  assign n19197 = n18983 & ~n19092;
  assign n19198 = ~n18977 & ~n19197;
  assign n19199 = ~n19196 & n19198;
  assign n19181 = n5942 & n10303;
  assign n19182 = x123 & n6186;
  assign n19183 = x124 & n5947;
  assign n19184 = ~n19182 & ~n19183;
  assign n19185 = x125 & n6406;
  assign n19186 = n19184 & ~n19185;
  assign n19187 = ~n19181 & n19186;
  assign n19188 = n19187 ^ x47;
  assign n19178 = n19070 ^ n19059;
  assign n19179 = n19071 & ~n19178;
  assign n19180 = n19179 ^ n19062;
  assign n19189 = n19188 ^ n19180;
  assign n19166 = n7395 & n8542;
  assign n19167 = x117 & n7650;
  assign n19168 = x118 & n7400;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = x119 & n7652;
  assign n19171 = n19169 & ~n19170;
  assign n19172 = ~n19166 & n19171;
  assign n19173 = n19172 ^ x53;
  assign n19156 = n7730 & n8171;
  assign n19157 = x114 & n8181;
  assign n19158 = x115 & n8174;
  assign n19159 = ~n19157 & ~n19158;
  assign n19160 = x116 & n8732;
  assign n19161 = n19159 & ~n19160;
  assign n19162 = ~n19156 & n19161;
  assign n19163 = n19162 ^ x56;
  assign n19153 = n19034 ^ n19003;
  assign n19154 = ~n19035 & n19153;
  assign n19155 = n19154 ^ n19003;
  assign n19164 = n19163 ^ n19155;
  assign n19143 = n6975 & n9002;
  assign n19144 = x111 & n9012;
  assign n19145 = x112 & n9005;
  assign n19146 = ~n19144 & ~n19145;
  assign n19147 = x113 & n9557;
  assign n19148 = n19146 & ~n19147;
  assign n19149 = ~n19143 & n19148;
  assign n19150 = n19149 ^ x59;
  assign n19140 = n19024 ^ n19013;
  assign n19141 = n19025 & ~n19140;
  assign n19142 = n19141 ^ n19016;
  assign n19151 = n19150 ^ n19142;
  assign n19131 = n6250 & n9878;
  assign n19132 = x109 & n9881;
  assign n19133 = x108 & n9888;
  assign n19134 = ~n19132 & ~n19133;
  assign n19135 = x110 & n10501;
  assign n19136 = n19134 & ~n19135;
  assign n19137 = ~n19131 & n19136;
  assign n19138 = n19137 ^ x62;
  assign n19123 = n5101 ^ x107;
  assign n19124 = x107 ^ x63;
  assign n19125 = n19124 ^ x107;
  assign n19126 = n19123 & n19125;
  assign n19127 = n19126 ^ x107;
  assign n19128 = ~n10177 & n19127;
  assign n19129 = n19128 ^ x107;
  assign n19120 = n18741 ^ x41;
  assign n19121 = ~n19012 & ~n19120;
  assign n19122 = n19121 ^ x41;
  assign n19130 = n19129 ^ n19122;
  assign n19139 = n19138 ^ n19130;
  assign n19152 = n19151 ^ n19139;
  assign n19165 = n19164 ^ n19152;
  assign n19174 = n19173 ^ n19165;
  assign n19117 = n19044 ^ n19000;
  assign n19118 = ~n19045 & n19117;
  assign n19119 = n19118 ^ n19000;
  assign n19175 = n19174 ^ n19119;
  assign n19114 = n19057 ^ n19046;
  assign n19115 = n19058 & ~n19114;
  assign n19116 = n19115 ^ n19049;
  assign n19176 = n19175 ^ n19116;
  assign n19106 = n6626 & n9387;
  assign n19107 = x120 & n6884;
  assign n19108 = x121 & n6630;
  assign n19109 = ~n19107 & ~n19108;
  assign n19110 = x122 & n6888;
  assign n19111 = n19109 & ~n19110;
  assign n19112 = ~n19106 & n19111;
  assign n19113 = n19112 ^ x50;
  assign n19177 = n19176 ^ n19113;
  assign n19190 = n19189 ^ n19177;
  assign n19103 = n19080 ^ n18997;
  assign n19104 = ~n19081 & n19103;
  assign n19105 = n19104 ^ n18997;
  assign n19191 = n19190 ^ n19105;
  assign n19097 = n5262 & ~n10281;
  assign n19098 = x127 & n5266;
  assign n19099 = x126 & n5488;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = ~n19097 & n19100;
  assign n19102 = n19101 ^ x44;
  assign n19192 = n19191 ^ n19102;
  assign n19094 = n19090 ^ n18994;
  assign n19095 = ~n19091 & n19094;
  assign n19096 = n19095 ^ n18994;
  assign n19193 = n19192 ^ n19096;
  assign n19200 = n19199 ^ n19193;
  assign n19294 = x127 & n5051;
  assign n19295 = ~x44 & ~n19294;
  assign n19296 = n19295 ^ x43;
  assign n19297 = n4848 & n11409;
  assign n19298 = n19297 ^ n19295;
  assign n19299 = ~n19295 & n19298;
  assign n19300 = n19299 ^ n19295;
  assign n19301 = x127 & n5487;
  assign n19302 = ~n19300 & ~n19301;
  assign n19303 = n19302 ^ n19299;
  assign n19304 = n19303 ^ n19295;
  assign n19305 = n19304 ^ n19297;
  assign n19306 = ~n19296 & n19305;
  assign n19307 = n19306 ^ x43;
  assign n19291 = n19180 ^ n19177;
  assign n19292 = n19189 & ~n19291;
  assign n19293 = n19292 ^ n19188;
  assign n19308 = n19307 ^ n19293;
  assign n19281 = n5942 & ~n10570;
  assign n19282 = x124 & n6186;
  assign n19283 = x126 & n6406;
  assign n19284 = ~n19282 & ~n19283;
  assign n19285 = x125 & n5947;
  assign n19286 = n19284 & ~n19285;
  assign n19287 = ~n19281 & n19286;
  assign n19288 = n19287 ^ x47;
  assign n19271 = n6626 & n9691;
  assign n19272 = x121 & n6884;
  assign n19273 = x122 & n6630;
  assign n19274 = ~n19272 & ~n19273;
  assign n19275 = x123 & n6888;
  assign n19276 = n19274 & ~n19275;
  assign n19277 = ~n19271 & n19276;
  assign n19278 = n19277 ^ x50;
  assign n19261 = n7395 & n8820;
  assign n19262 = x118 & n7650;
  assign n19263 = x119 & n7400;
  assign n19264 = ~n19262 & ~n19263;
  assign n19265 = x120 & n7652;
  assign n19266 = n19264 & ~n19265;
  assign n19267 = ~n19261 & n19266;
  assign n19268 = n19267 ^ x53;
  assign n19251 = n7987 & n8171;
  assign n19252 = x115 & n8181;
  assign n19253 = x116 & n8174;
  assign n19254 = ~n19252 & ~n19253;
  assign n19255 = x117 & n8732;
  assign n19256 = n19254 & ~n19255;
  assign n19257 = ~n19251 & n19256;
  assign n19258 = n19257 ^ x56;
  assign n19242 = n7220 & n9002;
  assign n19243 = x112 & n9012;
  assign n19244 = x113 & n9005;
  assign n19245 = ~n19243 & ~n19244;
  assign n19246 = x114 & n9557;
  assign n19247 = n19245 & ~n19246;
  assign n19248 = ~n19242 & n19247;
  assign n19249 = n19248 ^ x59;
  assign n19233 = n6478 & n9878;
  assign n19234 = x109 & n9888;
  assign n19235 = x111 & n10501;
  assign n19236 = ~n19234 & ~n19235;
  assign n19237 = x110 & n9881;
  assign n19238 = n19236 & ~n19237;
  assign n19239 = ~n19233 & n19238;
  assign n19222 = n5335 ^ x62;
  assign n19223 = n19222 ^ x63;
  assign n19224 = n19223 ^ n5335;
  assign n19225 = n5335 ^ x63;
  assign n19226 = n19225 ^ n5335;
  assign n19227 = n5335 ^ n5101;
  assign n19228 = n19227 ^ n5335;
  assign n19229 = n19226 & n19228;
  assign n19230 = n19229 ^ n5335;
  assign n19231 = ~n19224 & n19230;
  assign n19232 = n19231 ^ n19222;
  assign n19240 = n19239 ^ n19232;
  assign n19219 = n19138 ^ n19122;
  assign n19220 = ~n19130 & n19219;
  assign n19221 = n19220 ^ n19138;
  assign n19241 = n19240 ^ n19221;
  assign n19250 = n19249 ^ n19241;
  assign n19259 = n19258 ^ n19250;
  assign n19216 = n19142 ^ n19139;
  assign n19217 = n19151 & ~n19216;
  assign n19218 = n19217 ^ n19150;
  assign n19260 = n19259 ^ n19218;
  assign n19269 = n19268 ^ n19260;
  assign n19213 = n19155 ^ n19152;
  assign n19214 = n19164 & ~n19213;
  assign n19215 = n19214 ^ n19163;
  assign n19270 = n19269 ^ n19215;
  assign n19279 = n19278 ^ n19270;
  assign n19210 = n19165 ^ n19119;
  assign n19211 = n19174 & ~n19210;
  assign n19212 = n19211 ^ n19173;
  assign n19280 = n19279 ^ n19212;
  assign n19289 = n19288 ^ n19280;
  assign n19207 = n19175 ^ n19113;
  assign n19208 = n19176 & ~n19207;
  assign n19209 = n19208 ^ n19116;
  assign n19290 = n19289 ^ n19209;
  assign n19309 = n19308 ^ n19290;
  assign n19204 = n19190 ^ n19102;
  assign n19205 = n19191 & ~n19204;
  assign n19206 = n19205 ^ n19105;
  assign n19310 = n19309 ^ n19206;
  assign n19201 = n19199 ^ n19192;
  assign n19202 = n19193 & ~n19201;
  assign n19203 = n19202 ^ n19096;
  assign n19311 = n19310 ^ n19203;
  assign n19429 = n19206 & n19293;
  assign n19430 = n19307 ^ n19290;
  assign n19431 = ~n19206 & ~n19293;
  assign n19432 = n19431 ^ n19290;
  assign n19433 = n19430 & ~n19432;
  assign n19434 = n19433 ^ n19307;
  assign n19435 = ~n19429 & n19434;
  assign n19422 = n19290 & n19307;
  assign n19423 = n19293 ^ n19206;
  assign n19424 = ~n19290 & ~n19307;
  assign n19425 = n19424 ^ n19206;
  assign n19426 = n19423 & n19425;
  assign n19427 = n19426 ^ n19206;
  assign n19428 = ~n19422 & n19427;
  assign n19436 = n19435 ^ n19428;
  assign n19437 = n19203 & n19436;
  assign n19438 = n19437 ^ n19435;
  assign n19439 = n19431 ^ n19429;
  assign n19440 = n19433 ^ n19290;
  assign n19441 = n19439 & n19440;
  assign n19442 = n19441 ^ n19429;
  assign n19443 = ~n19438 & ~n19442;
  assign n19412 = n5942 & ~n10855;
  assign n19413 = x125 & n6186;
  assign n19414 = x126 & n5947;
  assign n19415 = ~n19413 & ~n19414;
  assign n19416 = x127 & n6406;
  assign n19417 = n19415 & ~n19416;
  assign n19418 = ~n19412 & n19417;
  assign n19419 = n19418 ^ x47;
  assign n19402 = n6626 & n9999;
  assign n19403 = x122 & n6884;
  assign n19404 = x123 & n6630;
  assign n19405 = ~n19403 & ~n19404;
  assign n19406 = x124 & n6888;
  assign n19407 = n19405 & ~n19406;
  assign n19408 = ~n19402 & n19407;
  assign n19409 = n19408 ^ x50;
  assign n19392 = n7395 & n9094;
  assign n19393 = x119 & n7650;
  assign n19394 = x120 & n7400;
  assign n19395 = ~n19393 & ~n19394;
  assign n19396 = x121 & n7652;
  assign n19397 = n19395 & ~n19396;
  assign n19398 = ~n19392 & n19397;
  assign n19399 = n19398 ^ x53;
  assign n19389 = n19260 ^ n19215;
  assign n19390 = ~n19269 & n19389;
  assign n19391 = n19390 ^ n19268;
  assign n19400 = n19399 ^ n19391;
  assign n19377 = n7481 & n9002;
  assign n19378 = x113 & n9012;
  assign n19379 = x114 & n9005;
  assign n19380 = ~n19378 & ~n19379;
  assign n19381 = x115 & n9557;
  assign n19382 = n19380 & ~n19381;
  assign n19383 = ~n19377 & n19382;
  assign n19384 = n19383 ^ x59;
  assign n19374 = n19249 ^ n19221;
  assign n19375 = n19241 & n19374;
  assign n19376 = n19375 ^ n19249;
  assign n19385 = n19384 ^ n19376;
  assign n19347 = ~x107 & x108;
  assign n19350 = n14116 & ~n19347;
  assign n19348 = x63 & n19347;
  assign n19349 = ~x62 & ~n19348;
  assign n19351 = n19350 ^ n19349;
  assign n19352 = x107 & ~x108;
  assign n19353 = n19352 ^ n19349;
  assign n19354 = n19349 ^ n19239;
  assign n19355 = ~n19349 & ~n19354;
  assign n19356 = n19355 ^ n19349;
  assign n19357 = ~n19353 & ~n19356;
  assign n19358 = n19357 ^ n19355;
  assign n19359 = n19358 ^ n19349;
  assign n19360 = n19359 ^ n19239;
  assign n19361 = n19351 & ~n19360;
  assign n19362 = n19361 ^ n19350;
  assign n19363 = n19352 ^ x62;
  assign n19364 = n19363 ^ n19352;
  assign n19365 = n19239 ^ x107;
  assign n19366 = ~n5101 & n19365;
  assign n19367 = n19366 ^ x107;
  assign n19368 = n19367 ^ n19352;
  assign n19369 = n19364 & ~n19368;
  assign n19370 = n19369 ^ n19352;
  assign n19371 = x63 & n19370;
  assign n19372 = ~n19362 & ~n19371;
  assign n19338 = n6728 & n9878;
  assign n19339 = x110 & n9888;
  assign n19340 = x112 & n10501;
  assign n19341 = ~n19339 & ~n19340;
  assign n19342 = x111 & n9881;
  assign n19343 = n19341 & ~n19342;
  assign n19344 = ~n19338 & n19343;
  assign n19345 = n19344 ^ x62;
  assign n19329 = n5554 ^ x109;
  assign n19330 = x109 ^ x63;
  assign n19331 = n19330 ^ x109;
  assign n19332 = n19329 & n19331;
  assign n19333 = n19332 ^ x109;
  assign n19334 = ~n10177 & n19333;
  assign n19335 = n19334 ^ x109;
  assign n19336 = n19335 ^ n19129;
  assign n19337 = n19336 ^ x44;
  assign n19346 = n19345 ^ n19337;
  assign n19373 = n19372 ^ n19346;
  assign n19386 = n19385 ^ n19373;
  assign n19321 = n8171 & n8265;
  assign n19322 = x116 & n8181;
  assign n19323 = x117 & n8174;
  assign n19324 = ~n19322 & ~n19323;
  assign n19325 = x118 & n8732;
  assign n19326 = n19324 & ~n19325;
  assign n19327 = ~n19321 & n19326;
  assign n19328 = n19327 ^ x56;
  assign n19387 = n19386 ^ n19328;
  assign n19318 = n19250 ^ n19218;
  assign n19319 = ~n19259 & n19318;
  assign n19320 = n19319 ^ n19258;
  assign n19388 = n19387 ^ n19320;
  assign n19401 = n19400 ^ n19388;
  assign n19410 = n19409 ^ n19401;
  assign n19315 = n19270 ^ n19212;
  assign n19316 = ~n19279 & n19315;
  assign n19317 = n19316 ^ n19278;
  assign n19411 = n19410 ^ n19317;
  assign n19420 = n19419 ^ n19411;
  assign n19312 = n19280 ^ n19209;
  assign n19313 = ~n19289 & n19312;
  assign n19314 = n19313 ^ n19288;
  assign n19421 = n19420 ^ n19314;
  assign n19444 = n19443 ^ n19421;
  assign n19528 = n19421 & ~n19429;
  assign n19529 = ~n19422 & ~n19528;
  assign n19530 = n19203 & n19529;
  assign n19531 = ~n19421 & ~n19434;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = n19421 & ~n19424;
  assign n19534 = n19206 ^ n19203;
  assign n19535 = n19423 & n19534;
  assign n19536 = n19535 ^ n19206;
  assign n19537 = ~n19533 & n19536;
  assign n19538 = n19532 & ~n19537;
  assign n19519 = n5942 & ~n10281;
  assign n19520 = x126 & n6186;
  assign n19521 = x127 & n5947;
  assign n19522 = ~n19520 & ~n19521;
  assign n19523 = ~n19519 & n19522;
  assign n19524 = n19523 ^ x47;
  assign n19509 = n6626 & n10303;
  assign n19510 = x123 & n6884;
  assign n19511 = x124 & n6630;
  assign n19512 = ~n19510 & ~n19511;
  assign n19513 = x125 & n6888;
  assign n19514 = n19512 & ~n19513;
  assign n19515 = ~n19509 & n19514;
  assign n19516 = n19515 ^ x50;
  assign n19499 = n7395 & n9387;
  assign n19500 = x120 & n7650;
  assign n19501 = x121 & n7400;
  assign n19502 = ~n19500 & ~n19501;
  assign n19503 = x122 & n7652;
  assign n19504 = n19502 & ~n19503;
  assign n19505 = ~n19499 & n19504;
  assign n19506 = n19505 ^ x53;
  assign n19489 = n8171 & n8542;
  assign n19490 = x117 & n8181;
  assign n19491 = x118 & n8174;
  assign n19492 = ~n19490 & ~n19491;
  assign n19493 = x119 & n8732;
  assign n19494 = n19492 & ~n19493;
  assign n19495 = ~n19489 & n19494;
  assign n19496 = n19495 ^ x56;
  assign n19479 = n7730 & n9002;
  assign n19480 = x114 & n9012;
  assign n19481 = x116 & n9557;
  assign n19482 = ~n19480 & ~n19481;
  assign n19483 = x115 & n9005;
  assign n19484 = n19482 & ~n19483;
  assign n19485 = ~n19479 & n19484;
  assign n19486 = n19485 ^ x59;
  assign n19469 = n6975 & n9878;
  assign n19470 = x111 & n9888;
  assign n19471 = x112 & n9881;
  assign n19472 = ~n19470 & ~n19471;
  assign n19473 = x113 & n10501;
  assign n19474 = n19472 & ~n19473;
  assign n19475 = ~n19469 & n19474;
  assign n19476 = n19475 ^ x62;
  assign n19466 = n19129 ^ x44;
  assign n19467 = ~n19336 & ~n19466;
  assign n19468 = n19467 ^ x44;
  assign n19477 = n19476 ^ n19468;
  assign n19463 = x110 & n10177;
  assign n19464 = x109 & n12123;
  assign n19465 = ~n19463 & ~n19464;
  assign n19478 = n19477 ^ n19465;
  assign n19487 = n19486 ^ n19478;
  assign n19460 = n19372 ^ n19345;
  assign n19461 = ~n19346 & ~n19460;
  assign n19462 = n19461 ^ n19372;
  assign n19488 = n19487 ^ n19462;
  assign n19497 = n19496 ^ n19488;
  assign n19457 = n19384 ^ n19373;
  assign n19458 = n19385 & n19457;
  assign n19459 = n19458 ^ n19376;
  assign n19498 = n19497 ^ n19459;
  assign n19507 = n19506 ^ n19498;
  assign n19454 = n19386 ^ n19320;
  assign n19455 = n19387 & ~n19454;
  assign n19456 = n19455 ^ n19320;
  assign n19508 = n19507 ^ n19456;
  assign n19517 = n19516 ^ n19508;
  assign n19451 = n19399 ^ n19388;
  assign n19452 = n19400 & n19451;
  assign n19453 = n19452 ^ n19391;
  assign n19518 = n19517 ^ n19453;
  assign n19525 = n19524 ^ n19518;
  assign n19448 = n19409 ^ n19317;
  assign n19449 = n19410 & n19448;
  assign n19450 = n19449 ^ n19317;
  assign n19526 = n19525 ^ n19450;
  assign n19445 = n19419 ^ n19314;
  assign n19446 = n19420 & n19445;
  assign n19447 = n19446 ^ n19314;
  assign n19527 = n19526 ^ n19447;
  assign n19539 = n19538 ^ n19527;
  assign n19629 = ~n19518 & ~n19524;
  assign n19630 = n19447 & n19450;
  assign n19642 = n19629 & ~n19630;
  assign n19632 = ~n19447 & ~n19450;
  assign n19634 = n19518 & n19524;
  assign n19643 = n19632 & ~n19634;
  assign n19644 = ~n19642 & ~n19643;
  assign n19631 = n19630 ^ n19629;
  assign n19633 = n19632 ^ n19631;
  assign n19635 = n19634 ^ n19633;
  assign n19636 = n19632 ^ n19629;
  assign n19637 = n19634 ^ n19632;
  assign n19638 = ~n19636 & n19637;
  assign n19639 = ~n19635 & n19638;
  assign n19640 = n19639 ^ n19635;
  assign n19641 = ~n19538 & n19640;
  assign n19645 = n19644 ^ n19641;
  assign n19646 = n19632 ^ n19630;
  assign n19647 = n19630 ^ n19518;
  assign n19648 = n19647 ^ n19630;
  assign n19649 = n19646 & ~n19648;
  assign n19650 = n19649 ^ n19630;
  assign n19651 = ~n19525 & n19650;
  assign n19652 = n19645 & ~n19651;
  assign n19617 = n6626 & ~n10570;
  assign n19618 = x124 & n6884;
  assign n19619 = x126 & n6888;
  assign n19620 = ~n19618 & ~n19619;
  assign n19621 = x125 & n6630;
  assign n19622 = n19620 & ~n19621;
  assign n19623 = ~n19617 & n19622;
  assign n19624 = n19623 ^ x50;
  assign n19607 = n7395 & n9691;
  assign n19608 = x121 & n7650;
  assign n19609 = x122 & n7400;
  assign n19610 = ~n19608 & ~n19609;
  assign n19611 = x123 & n7652;
  assign n19612 = n19610 & ~n19611;
  assign n19613 = ~n19607 & n19612;
  assign n19614 = n19613 ^ x53;
  assign n19597 = n8171 & n8820;
  assign n19598 = x118 & n8181;
  assign n19599 = x119 & n8174;
  assign n19600 = ~n19598 & ~n19599;
  assign n19601 = x120 & n8732;
  assign n19602 = n19600 & ~n19601;
  assign n19603 = ~n19597 & n19602;
  assign n19604 = n19603 ^ x56;
  assign n19594 = n19478 ^ n19462;
  assign n19595 = ~n19487 & ~n19594;
  assign n19596 = n19595 ^ n19486;
  assign n19605 = n19604 ^ n19596;
  assign n19584 = n7987 & n9002;
  assign n19585 = x115 & n9012;
  assign n19586 = x117 & n9557;
  assign n19587 = ~n19585 & ~n19586;
  assign n19588 = x116 & n9005;
  assign n19589 = n19587 & ~n19588;
  assign n19590 = ~n19584 & n19589;
  assign n19591 = n19590 ^ x59;
  assign n19576 = n7220 & n9878;
  assign n19577 = x112 & n9888;
  assign n19578 = x113 & n9881;
  assign n19579 = ~n19577 & ~n19578;
  assign n19580 = x114 & n10501;
  assign n19581 = n19579 & ~n19580;
  assign n19582 = ~n19576 & n19581;
  assign n19583 = n19582 ^ x62;
  assign n19592 = n19591 ^ n19583;
  assign n19572 = n19468 ^ n19465;
  assign n19573 = n19477 & n19572;
  assign n19574 = n19573 ^ n19476;
  assign n19563 = x111 ^ x110;
  assign n19564 = n19563 ^ x63;
  assign n19565 = n19564 ^ n19563;
  assign n19566 = n19563 ^ n6249;
  assign n19567 = n19566 ^ n19563;
  assign n19568 = n19565 & n19567;
  assign n19569 = n19568 ^ n19563;
  assign n19570 = ~n10177 & n19569;
  assign n19571 = n19570 ^ n19563;
  assign n19575 = n19574 ^ n19571;
  assign n19593 = n19592 ^ n19575;
  assign n19606 = n19605 ^ n19593;
  assign n19615 = n19614 ^ n19606;
  assign n19560 = n19488 ^ n19459;
  assign n19561 = n19497 & ~n19560;
  assign n19562 = n19561 ^ n19496;
  assign n19616 = n19615 ^ n19562;
  assign n19625 = n19624 ^ n19616;
  assign n19557 = n19498 ^ n19456;
  assign n19558 = n19507 & ~n19557;
  assign n19559 = n19558 ^ n19506;
  assign n19626 = n19625 ^ n19559;
  assign n19543 = x127 & n5709;
  assign n19544 = ~x47 & ~n19543;
  assign n19545 = n19544 ^ x46;
  assign n19546 = n5481 & n11409;
  assign n19547 = n19546 ^ n19544;
  assign n19548 = ~n19544 & n19547;
  assign n19549 = n19548 ^ n19544;
  assign n19550 = x127 & n6185;
  assign n19551 = ~n19549 & ~n19550;
  assign n19552 = n19551 ^ n19548;
  assign n19553 = n19552 ^ n19544;
  assign n19554 = n19553 ^ n19546;
  assign n19555 = ~n19545 & n19554;
  assign n19556 = n19555 ^ x46;
  assign n19627 = n19626 ^ n19556;
  assign n19540 = n19508 ^ n19453;
  assign n19541 = n19517 & ~n19540;
  assign n19542 = n19541 ^ n19516;
  assign n19628 = n19627 ^ n19542;
  assign n19653 = n19652 ^ n19628;
  assign n19749 = n19628 & ~n19643;
  assign n19750 = n19538 & ~n19749;
  assign n19751 = ~n19628 & ~n19630;
  assign n19752 = ~n19629 & ~n19751;
  assign n19753 = ~n19750 & n19752;
  assign n19754 = ~n19628 & ~n19634;
  assign n19755 = n19538 ^ n19447;
  assign n19756 = n19450 ^ n19447;
  assign n19757 = ~n19755 & n19756;
  assign n19758 = n19757 ^ n19447;
  assign n19759 = ~n19754 & n19758;
  assign n19760 = ~n19753 & ~n19759;
  assign n19744 = n19626 ^ n19542;
  assign n19745 = n19627 & n19744;
  assign n19746 = n19745 ^ n19556;
  assign n19741 = n19616 ^ n19559;
  assign n19742 = ~n19625 & n19741;
  assign n19743 = n19742 ^ n19624;
  assign n19747 = n19746 ^ n19743;
  assign n19732 = n6626 & ~n10855;
  assign n19733 = x125 & n6884;
  assign n19734 = x126 & n6630;
  assign n19735 = ~n19733 & ~n19734;
  assign n19736 = x127 & n6888;
  assign n19737 = n19735 & ~n19736;
  assign n19738 = ~n19732 & n19737;
  assign n19739 = n19738 ^ x50;
  assign n19722 = n7395 & n9999;
  assign n19723 = x122 & n7650;
  assign n19724 = x124 & n7652;
  assign n19725 = ~n19723 & ~n19724;
  assign n19726 = x123 & n7400;
  assign n19727 = n19725 & ~n19726;
  assign n19728 = ~n19722 & n19727;
  assign n19729 = n19728 ^ x53;
  assign n19710 = n8265 & n9002;
  assign n19711 = x116 & n9012;
  assign n19712 = x118 & n9557;
  assign n19713 = ~n19711 & ~n19712;
  assign n19714 = x117 & n9005;
  assign n19715 = n19713 & ~n19714;
  assign n19716 = ~n19710 & n19715;
  assign n19717 = n19716 ^ x59;
  assign n19707 = n19583 ^ n19575;
  assign n19708 = n19592 & n19707;
  assign n19709 = n19708 ^ n19591;
  assign n19718 = n19717 ^ n19709;
  assign n19686 = n19464 ^ x111;
  assign n19687 = n19686 ^ n19464;
  assign n19688 = n19464 ^ n10177;
  assign n19689 = n19688 ^ n19464;
  assign n19690 = ~n19687 & n19689;
  assign n19691 = n19690 ^ n19464;
  assign n19692 = x110 & n19691;
  assign n19693 = n19692 ^ n19464;
  assign n19694 = n19574 & ~n19693;
  assign n19695 = n10177 ^ x110;
  assign n19696 = n19563 ^ x111;
  assign n19697 = n19696 ^ n19695;
  assign n19698 = ~x109 & ~n19330;
  assign n19699 = n19698 ^ x111;
  assign n19700 = n19699 ^ x109;
  assign n19701 = n19697 & ~n19700;
  assign n19702 = n19701 ^ n19698;
  assign n19703 = n19702 ^ x109;
  assign n19704 = n19695 & ~n19703;
  assign n19705 = ~n19694 & ~n19704;
  assign n19677 = n7481 & n9878;
  assign n19678 = x113 & n9888;
  assign n19679 = x114 & n9881;
  assign n19680 = ~n19678 & ~n19679;
  assign n19681 = x115 & n10501;
  assign n19682 = n19680 & ~n19681;
  assign n19683 = ~n19677 & n19682;
  assign n19684 = n19683 ^ x62;
  assign n19668 = n19563 ^ n6232;
  assign n19669 = n19668 ^ n6232;
  assign n19670 = n6232 ^ x63;
  assign n19671 = n19670 ^ n6232;
  assign n19672 = n19669 & n19671;
  assign n19673 = n19672 ^ n6232;
  assign n19674 = ~n10177 & n19673;
  assign n19675 = n19674 ^ n6232;
  assign n19676 = n19675 ^ x47;
  assign n19685 = n19684 ^ n19676;
  assign n19706 = n19705 ^ n19685;
  assign n19719 = n19718 ^ n19706;
  assign n19660 = n8171 & n9094;
  assign n19661 = x119 & n8181;
  assign n19662 = x121 & n8732;
  assign n19663 = ~n19661 & ~n19662;
  assign n19664 = x120 & n8174;
  assign n19665 = n19663 & ~n19664;
  assign n19666 = ~n19660 & n19665;
  assign n19667 = n19666 ^ x56;
  assign n19720 = n19719 ^ n19667;
  assign n19657 = n19604 ^ n19593;
  assign n19658 = n19605 & n19657;
  assign n19659 = n19658 ^ n19596;
  assign n19721 = n19720 ^ n19659;
  assign n19730 = n19729 ^ n19721;
  assign n19654 = n19606 ^ n19562;
  assign n19655 = ~n19615 & n19654;
  assign n19656 = n19655 ^ n19614;
  assign n19731 = n19730 ^ n19656;
  assign n19740 = n19739 ^ n19731;
  assign n19748 = n19747 ^ n19740;
  assign n19761 = n19760 ^ n19748;
  assign n19838 = n19731 & ~n19739;
  assign n19839 = ~n19760 & ~n19838;
  assign n19840 = ~n19731 & n19739;
  assign n19841 = n19840 ^ n19743;
  assign n19842 = ~n19747 & ~n19841;
  assign n19843 = n19842 ^ n19746;
  assign n19844 = n19839 & ~n19843;
  assign n19845 = n19743 & ~n19746;
  assign n19846 = n19838 & ~n19845;
  assign n19847 = ~n19743 & n19746;
  assign n19848 = ~n19840 & n19847;
  assign n19849 = ~n19846 & ~n19848;
  assign n19850 = n19760 & ~n19849;
  assign n19851 = n19847 ^ n19845;
  assign n19852 = n19845 ^ n19731;
  assign n19853 = n19852 ^ n19845;
  assign n19854 = n19851 & n19853;
  assign n19855 = n19854 ^ n19845;
  assign n19856 = n19740 & n19855;
  assign n19857 = ~n19850 & ~n19856;
  assign n19858 = ~n19844 & n19857;
  assign n19826 = n7395 & n10303;
  assign n19827 = x123 & n7650;
  assign n19828 = x125 & n7652;
  assign n19829 = ~n19827 & ~n19828;
  assign n19830 = x124 & n7400;
  assign n19831 = n19829 & ~n19830;
  assign n19832 = ~n19826 & n19831;
  assign n19833 = n19832 ^ x53;
  assign n19823 = n19667 ^ n19659;
  assign n19824 = ~n19720 & ~n19823;
  assign n19825 = n19824 ^ n19719;
  assign n19834 = n19833 ^ n19825;
  assign n19813 = n8171 & n9387;
  assign n19814 = x120 & n8181;
  assign n19815 = x121 & n8174;
  assign n19816 = ~n19814 & ~n19815;
  assign n19817 = x122 & n8732;
  assign n19818 = n19816 & ~n19817;
  assign n19819 = ~n19813 & n19818;
  assign n19820 = n19819 ^ x56;
  assign n19810 = n19717 ^ n19706;
  assign n19811 = n19718 & n19810;
  assign n19812 = n19811 ^ n19709;
  assign n19821 = n19820 ^ n19812;
  assign n19800 = n8542 & n9002;
  assign n19801 = x118 & n9005;
  assign n19802 = x117 & n9012;
  assign n19803 = ~n19801 & ~n19802;
  assign n19804 = x119 & n9557;
  assign n19805 = n19803 & ~n19804;
  assign n19806 = ~n19800 & n19805;
  assign n19807 = n19806 ^ x59;
  assign n19791 = n7730 & n9878;
  assign n19792 = x114 & n9888;
  assign n19793 = x115 & n9881;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = x116 & n10501;
  assign n19796 = n19794 & ~n19795;
  assign n19797 = ~n19791 & n19796;
  assign n19798 = n19797 ^ x62;
  assign n19782 = x111 ^ x47;
  assign n19783 = x112 ^ x110;
  assign n19784 = ~n12123 & n19783;
  assign n19785 = n19784 ^ x110;
  assign n19786 = n19785 ^ x111;
  assign n19787 = ~n19782 & n19786;
  assign n19788 = n19787 ^ x111;
  assign n19789 = ~n12893 & n19788;
  assign n19774 = x113 ^ x112;
  assign n19775 = n19774 ^ x113;
  assign n19776 = x113 ^ x63;
  assign n19777 = n19776 ^ x113;
  assign n19778 = n19775 & n19777;
  assign n19779 = n19778 ^ x113;
  assign n19780 = ~n10177 & n19779;
  assign n19781 = n19780 ^ x113;
  assign n19790 = n19789 ^ n19781;
  assign n19799 = n19798 ^ n19790;
  assign n19808 = n19807 ^ n19799;
  assign n19771 = n19705 ^ n19684;
  assign n19772 = ~n19685 & ~n19771;
  assign n19773 = n19772 ^ n19705;
  assign n19809 = n19808 ^ n19773;
  assign n19822 = n19821 ^ n19809;
  assign n19835 = n19834 ^ n19822;
  assign n19768 = n19729 ^ n19656;
  assign n19769 = n19730 & n19768;
  assign n19770 = n19769 ^ n19656;
  assign n19836 = n19835 ^ n19770;
  assign n19762 = n6626 & ~n10281;
  assign n19763 = x127 & n6630;
  assign n19764 = x126 & n6884;
  assign n19765 = ~n19763 & ~n19764;
  assign n19766 = ~n19762 & n19765;
  assign n19767 = n19766 ^ x50;
  assign n19837 = n19836 ^ n19767;
  assign n19859 = n19858 ^ n19837;
  assign n19941 = ~n19837 & ~n19847;
  assign n19942 = ~n19840 & ~n19941;
  assign n19943 = ~n19839 & n19942;
  assign n19944 = ~n19837 & ~n19838;
  assign n19945 = ~n19845 & ~n19944;
  assign n19946 = n19760 & n19945;
  assign n19947 = n19837 & n19843;
  assign n19948 = ~n19946 & ~n19947;
  assign n19949 = ~n19943 & n19948;
  assign n19929 = n7395 & ~n10570;
  assign n19930 = x124 & n7650;
  assign n19931 = x125 & n7400;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = x126 & n7652;
  assign n19934 = n19932 & ~n19933;
  assign n19935 = ~n19929 & n19934;
  assign n19936 = n19935 ^ x53;
  assign n19926 = n19820 ^ n19809;
  assign n19927 = n19821 & ~n19926;
  assign n19928 = n19927 ^ n19812;
  assign n19937 = n19936 ^ n19928;
  assign n19916 = n8171 & n9691;
  assign n19917 = x121 & n8181;
  assign n19918 = x123 & n8732;
  assign n19919 = ~n19917 & ~n19918;
  assign n19920 = x122 & n8174;
  assign n19921 = n19919 & ~n19920;
  assign n19922 = ~n19916 & n19921;
  assign n19923 = n19922 ^ x56;
  assign n19907 = n8820 & n9002;
  assign n19908 = x118 & n9012;
  assign n19909 = x119 & n9005;
  assign n19910 = ~n19908 & ~n19909;
  assign n19911 = x120 & n9557;
  assign n19912 = n19910 & ~n19911;
  assign n19913 = ~n19907 & n19912;
  assign n19914 = n19913 ^ x59;
  assign n19894 = n6709 ^ x62;
  assign n19895 = n19894 ^ x63;
  assign n19896 = n19895 ^ n6709;
  assign n19897 = n19774 ^ n6709;
  assign n19898 = n19897 ^ n6709;
  assign n19899 = n6709 ^ x63;
  assign n19900 = n19899 ^ n6709;
  assign n19901 = n19898 & n19900;
  assign n19902 = n19901 ^ n6709;
  assign n19903 = ~n19896 & n19902;
  assign n19904 = n19903 ^ n19894;
  assign n19887 = n7987 & n9878;
  assign n19888 = x115 & n9888;
  assign n19889 = x117 & n10501;
  assign n19890 = ~n19888 & ~n19889;
  assign n19891 = x116 & n9881;
  assign n19892 = n19890 & ~n19891;
  assign n19893 = ~n19887 & n19892;
  assign n19905 = n19904 ^ n19893;
  assign n19884 = n19798 ^ n19789;
  assign n19885 = n19790 & ~n19884;
  assign n19886 = n19885 ^ n19798;
  assign n19906 = n19905 ^ n19886;
  assign n19915 = n19914 ^ n19906;
  assign n19924 = n19923 ^ n19915;
  assign n19881 = n19807 ^ n19773;
  assign n19882 = n19808 & ~n19881;
  assign n19883 = n19882 ^ n19773;
  assign n19925 = n19924 ^ n19883;
  assign n19938 = n19937 ^ n19925;
  assign n19878 = n19835 ^ n19767;
  assign n19879 = ~n19836 & n19878;
  assign n19880 = n19879 ^ n19770;
  assign n19939 = n19938 ^ n19880;
  assign n19863 = x127 & n6411;
  assign n19864 = ~x50 & ~n19863;
  assign n19865 = n19864 ^ x49;
  assign n19866 = n6191 & n11409;
  assign n19867 = n19866 ^ n19864;
  assign n19868 = ~n19864 & n19867;
  assign n19869 = n19868 ^ n19864;
  assign n19870 = x127 & n6883;
  assign n19871 = ~n19869 & ~n19870;
  assign n19872 = n19871 ^ n19868;
  assign n19873 = n19872 ^ n19864;
  assign n19874 = n19873 ^ n19866;
  assign n19875 = ~n19865 & n19874;
  assign n19876 = n19875 ^ x49;
  assign n19860 = n19825 ^ n19822;
  assign n19861 = ~n19834 & n19860;
  assign n19862 = n19861 ^ n19833;
  assign n19877 = n19876 ^ n19862;
  assign n19940 = n19939 ^ n19877;
  assign n19950 = n19949 ^ n19940;
  assign n20030 = n19862 & ~n19876;
  assign n20031 = ~n19949 & ~n20030;
  assign n20032 = ~n19862 & n19876;
  assign n20033 = n20032 ^ n19938;
  assign n20034 = n19939 & n20033;
  assign n20035 = n20034 ^ n19880;
  assign n20036 = n20031 & ~n20035;
  assign n20037 = ~n19880 & ~n19938;
  assign n20038 = n20030 & ~n20037;
  assign n20039 = n19880 & n19938;
  assign n20040 = ~n20032 & n20039;
  assign n20041 = ~n20038 & ~n20040;
  assign n20042 = n19949 & ~n20041;
  assign n20043 = n20039 ^ n20037;
  assign n20044 = n20039 ^ n19862;
  assign n20045 = n20044 ^ n20039;
  assign n20046 = n20043 & ~n20045;
  assign n20047 = n20046 ^ n20039;
  assign n20048 = n19877 & n20047;
  assign n20049 = ~n20042 & ~n20048;
  assign n20050 = ~n20036 & n20049;
  assign n20020 = n7395 & ~n10855;
  assign n20021 = x125 & n7650;
  assign n20022 = x126 & n7400;
  assign n20023 = ~n20021 & ~n20022;
  assign n20024 = x127 & n7652;
  assign n20025 = n20023 & ~n20024;
  assign n20026 = ~n20020 & n20025;
  assign n20027 = n20026 ^ x53;
  assign n20010 = n8171 & n9999;
  assign n20011 = x122 & n8181;
  assign n20012 = x123 & n8174;
  assign n20013 = ~n20011 & ~n20012;
  assign n20014 = x124 & n8732;
  assign n20015 = n20013 & ~n20014;
  assign n20016 = ~n20010 & n20015;
  assign n20017 = n20016 ^ x56;
  assign n20000 = n9002 & n9094;
  assign n20001 = x120 & n9005;
  assign n20002 = x119 & n9012;
  assign n20003 = ~n20001 & ~n20002;
  assign n20004 = x121 & n9557;
  assign n20005 = n20003 & ~n20004;
  assign n20006 = ~n20000 & n20005;
  assign n20007 = n20006 ^ x59;
  assign n19997 = n19914 ^ n19886;
  assign n19998 = n19906 & n19997;
  assign n19999 = n19998 ^ n19914;
  assign n20008 = n20007 ^ n19999;
  assign n19976 = ~x113 & x114;
  assign n19977 = x63 & n19976;
  assign n19978 = ~x62 & ~n19977;
  assign n19979 = n19893 & n19978;
  assign n19980 = n19893 ^ x114;
  assign n19981 = ~n6709 & n19980;
  assign n19982 = n19981 ^ x114;
  assign n19983 = n14116 & ~n19982;
  assign n19984 = ~n19979 & ~n19983;
  assign n19985 = x113 & ~x114;
  assign n19986 = n19985 ^ x62;
  assign n19987 = n19986 ^ n19985;
  assign n19988 = n19893 ^ x113;
  assign n19989 = ~n19774 & n19988;
  assign n19990 = n19989 ^ x113;
  assign n19991 = n19990 ^ n19985;
  assign n19992 = n19987 & ~n19991;
  assign n19993 = n19992 ^ n19985;
  assign n19994 = x63 & n19993;
  assign n19995 = n19984 & ~n19994;
  assign n19967 = n8265 & n9878;
  assign n19968 = x116 & n9888;
  assign n19969 = x118 & n10501;
  assign n19970 = ~n19968 & ~n19969;
  assign n19971 = x117 & n9881;
  assign n19972 = n19970 & ~n19971;
  assign n19973 = ~n19967 & n19972;
  assign n19974 = n19973 ^ x62;
  assign n19957 = x115 ^ x114;
  assign n19958 = n19957 ^ x115;
  assign n19959 = x115 ^ x63;
  assign n19960 = n19959 ^ x115;
  assign n19961 = n19958 & n19960;
  assign n19962 = n19961 ^ x115;
  assign n19963 = ~n10177 & n19962;
  assign n19964 = n19963 ^ x115;
  assign n19965 = n19964 ^ x50;
  assign n19966 = n19965 ^ n19781;
  assign n19975 = n19974 ^ n19966;
  assign n19996 = n19995 ^ n19975;
  assign n20009 = n20008 ^ n19996;
  assign n20018 = n20017 ^ n20009;
  assign n19954 = n19915 ^ n19883;
  assign n19955 = ~n19924 & ~n19954;
  assign n19956 = n19955 ^ n19923;
  assign n20019 = n20018 ^ n19956;
  assign n20028 = n20027 ^ n20019;
  assign n19951 = n19928 ^ n19925;
  assign n19952 = n19937 & ~n19951;
  assign n19953 = n19952 ^ n19936;
  assign n20029 = n20028 ^ n19953;
  assign n20051 = n20050 ^ n20029;
  assign n20110 = n20029 & ~n20039;
  assign n20111 = ~n20032 & ~n20110;
  assign n20112 = ~n20031 & n20111;
  assign n20113 = n20029 & ~n20030;
  assign n20114 = ~n20037 & ~n20113;
  assign n20115 = n19949 & n20114;
  assign n20116 = ~n20029 & n20035;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = ~n20112 & n20117;
  assign n20097 = n8171 & n10303;
  assign n20098 = x123 & n8181;
  assign n20099 = x124 & n8174;
  assign n20100 = ~n20098 & ~n20099;
  assign n20101 = x125 & n8732;
  assign n20102 = n20100 & ~n20101;
  assign n20103 = ~n20097 & n20102;
  assign n20104 = n20103 ^ x56;
  assign n20094 = n20007 ^ n19996;
  assign n20095 = n20008 & n20094;
  assign n20096 = n20095 ^ n19999;
  assign n20105 = n20104 ^ n20096;
  assign n20084 = n9002 & n9387;
  assign n20085 = x120 & n9012;
  assign n20086 = x121 & n9005;
  assign n20087 = ~n20085 & ~n20086;
  assign n20088 = x122 & n9557;
  assign n20089 = n20087 & ~n20088;
  assign n20090 = ~n20084 & n20089;
  assign n20091 = n20090 ^ x59;
  assign n20074 = n8542 & n9878;
  assign n20075 = x117 & n9888;
  assign n20076 = x118 & n9881;
  assign n20077 = ~n20075 & ~n20076;
  assign n20078 = x119 & n10501;
  assign n20079 = n20077 & ~n20078;
  assign n20080 = ~n20074 & n20079;
  assign n20081 = n20080 ^ x62;
  assign n20070 = n19781 ^ x50;
  assign n20071 = n19964 ^ n19781;
  assign n20072 = ~n20070 & ~n20071;
  assign n20073 = n20072 ^ x50;
  assign n20082 = n20081 ^ n20073;
  assign n20067 = x115 & n12123;
  assign n20068 = x116 & n10177;
  assign n20069 = ~n20067 & ~n20068;
  assign n20083 = n20082 ^ n20069;
  assign n20092 = n20091 ^ n20083;
  assign n20064 = n19995 ^ n19974;
  assign n20065 = ~n19975 & ~n20064;
  assign n20066 = n20065 ^ n19995;
  assign n20093 = n20092 ^ n20066;
  assign n20106 = n20105 ^ n20093;
  assign n20061 = n20017 ^ n19956;
  assign n20062 = n20018 & n20061;
  assign n20063 = n20062 ^ n19956;
  assign n20107 = n20106 ^ n20063;
  assign n20055 = n7395 & ~n10281;
  assign n20056 = x127 & n7400;
  assign n20057 = x126 & n7650;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = ~n20055 & n20058;
  assign n20060 = n20059 ^ x53;
  assign n20108 = n20107 ^ n20060;
  assign n20052 = n20027 ^ n19953;
  assign n20053 = n20028 & n20052;
  assign n20054 = n20053 ^ n19953;
  assign n20109 = n20108 ^ n20054;
  assign n20119 = n20118 ^ n20109;
  assign n20198 = n20118 ^ n20108;
  assign n20199 = n20109 & n20198;
  assign n20200 = n20199 ^ n20054;
  assign n20186 = n8171 & ~n10570;
  assign n20187 = x124 & n8181;
  assign n20188 = x126 & n8732;
  assign n20189 = ~n20187 & ~n20188;
  assign n20190 = x125 & n8174;
  assign n20191 = n20189 & ~n20190;
  assign n20192 = ~n20186 & n20191;
  assign n20193 = n20192 ^ x56;
  assign n20175 = n9002 & n9691;
  assign n20176 = x121 & n9012;
  assign n20177 = x122 & n9005;
  assign n20178 = ~n20176 & ~n20177;
  assign n20179 = x123 & n9557;
  assign n20180 = n20178 & ~n20179;
  assign n20181 = ~n20175 & n20180;
  assign n20182 = n20181 ^ x59;
  assign n20167 = n8820 & n9878;
  assign n20168 = x118 & n9888;
  assign n20169 = x119 & n9881;
  assign n20170 = ~n20168 & ~n20169;
  assign n20171 = x120 & n10501;
  assign n20172 = n20170 & ~n20171;
  assign n20173 = ~n20167 & n20172;
  assign n20174 = n20173 ^ x62;
  assign n20183 = n20182 ^ n20174;
  assign n20146 = n20067 ^ x117;
  assign n20147 = n20146 ^ n20067;
  assign n20148 = n20067 ^ n10177;
  assign n20149 = n20148 ^ n20067;
  assign n20150 = ~n20147 & n20149;
  assign n20151 = n20150 ^ n20067;
  assign n20152 = x116 & n20151;
  assign n20153 = n20152 ^ n20067;
  assign n20154 = n10177 ^ x116;
  assign n20155 = x117 ^ x116;
  assign n20156 = n20155 ^ x117;
  assign n20157 = n20156 ^ n20154;
  assign n20158 = ~x115 & ~n19959;
  assign n20159 = n20158 ^ x117;
  assign n20160 = n20159 ^ x115;
  assign n20161 = n20157 & ~n20160;
  assign n20162 = n20161 ^ n20158;
  assign n20163 = n20162 ^ x115;
  assign n20164 = n20154 & ~n20163;
  assign n20165 = ~n20153 & ~n20164;
  assign n20143 = n20073 ^ n20069;
  assign n20144 = n20082 & n20143;
  assign n20145 = n20144 ^ n20081;
  assign n20166 = n20165 ^ n20145;
  assign n20184 = n20183 ^ n20166;
  assign n20140 = n20083 ^ n20066;
  assign n20141 = ~n20092 & ~n20140;
  assign n20142 = n20141 ^ n20091;
  assign n20185 = n20184 ^ n20142;
  assign n20194 = n20193 ^ n20185;
  assign n20126 = x127 & n7130;
  assign n20127 = ~x53 & ~n20126;
  assign n20128 = n20127 ^ x52;
  assign n20129 = n6878 & n11409;
  assign n20130 = n20129 ^ n20127;
  assign n20131 = ~n20127 & n20130;
  assign n20132 = n20131 ^ n20127;
  assign n20133 = x127 & n7649;
  assign n20134 = ~n20132 & ~n20133;
  assign n20135 = n20134 ^ n20131;
  assign n20136 = n20135 ^ n20127;
  assign n20137 = n20136 ^ n20129;
  assign n20138 = ~n20128 & n20137;
  assign n20139 = n20138 ^ x52;
  assign n20195 = n20194 ^ n20139;
  assign n20123 = n20096 ^ n20093;
  assign n20124 = n20105 & ~n20123;
  assign n20125 = n20124 ^ n20104;
  assign n20196 = n20195 ^ n20125;
  assign n20120 = n20106 ^ n20060;
  assign n20121 = n20107 & ~n20120;
  assign n20122 = n20121 ^ n20063;
  assign n20197 = n20196 ^ n20122;
  assign n20201 = n20200 ^ n20197;
  assign n20251 = n20194 ^ n20125;
  assign n20252 = ~n20195 & ~n20251;
  assign n20253 = n20252 ^ n20139;
  assign n20248 = n20193 ^ n20142;
  assign n20249 = ~n20185 & n20248;
  assign n20250 = n20249 ^ n20193;
  assign n20254 = n20253 ^ n20250;
  assign n20237 = n9002 & n9999;
  assign n20238 = x122 & n9012;
  assign n20239 = x123 & n9005;
  assign n20240 = ~n20238 & ~n20239;
  assign n20241 = x124 & n9557;
  assign n20242 = n20240 & ~n20241;
  assign n20243 = ~n20237 & n20242;
  assign n20244 = n20243 ^ x59;
  assign n20234 = n20174 ^ n20166;
  assign n20235 = n20183 & ~n20234;
  assign n20236 = n20235 ^ n20182;
  assign n20245 = n20244 ^ n20236;
  assign n20224 = n9094 & n9878;
  assign n20225 = x119 & n9888;
  assign n20226 = x120 & n9881;
  assign n20227 = ~n20225 & ~n20226;
  assign n20228 = x121 & n10501;
  assign n20229 = n20227 & ~n20228;
  assign n20230 = ~n20224 & n20229;
  assign n20231 = n20230 ^ x62;
  assign n20215 = n20155 ^ n7713;
  assign n20216 = n20215 ^ n7713;
  assign n20217 = n7713 ^ x63;
  assign n20218 = n20217 ^ n7713;
  assign n20219 = n20216 & n20218;
  assign n20220 = n20219 ^ n7713;
  assign n20221 = ~n10177 & n20220;
  assign n20222 = n20221 ^ n7713;
  assign n20223 = n20222 ^ x53;
  assign n20232 = n20231 ^ n20223;
  assign n20213 = n20145 & n20165;
  assign n20214 = n20213 ^ n20164;
  assign n20233 = n20232 ^ n20214;
  assign n20246 = n20245 ^ n20233;
  assign n20205 = n8171 & ~n10855;
  assign n20206 = x125 & n8181;
  assign n20207 = x127 & n8732;
  assign n20208 = ~n20206 & ~n20207;
  assign n20209 = x126 & n8174;
  assign n20210 = n20208 & ~n20209;
  assign n20211 = ~n20205 & n20210;
  assign n20212 = n20211 ^ x56;
  assign n20247 = n20246 ^ n20212;
  assign n20255 = n20254 ^ n20247;
  assign n20202 = n20200 ^ n20196;
  assign n20203 = ~n20197 & n20202;
  assign n20204 = n20203 ^ n20122;
  assign n20256 = n20255 ^ n20204;
  assign n20306 = ~n20212 & ~n20246;
  assign n20307 = n20204 & ~n20306;
  assign n20308 = ~n20250 & n20253;
  assign n20309 = n20212 & n20246;
  assign n20310 = ~n20308 & n20309;
  assign n20311 = n20250 & ~n20253;
  assign n20312 = ~n20310 & ~n20311;
  assign n20313 = n20307 & ~n20312;
  assign n20314 = n20306 & ~n20311;
  assign n20315 = ~n20308 & ~n20314;
  assign n20316 = ~n20309 & ~n20315;
  assign n20317 = ~n20204 & n20316;
  assign n20318 = ~n20310 & ~n20314;
  assign n20319 = n20254 & ~n20318;
  assign n20320 = ~n20317 & ~n20319;
  assign n20321 = ~n20313 & n20320;
  assign n20294 = n9002 & n10303;
  assign n20295 = x123 & n9012;
  assign n20296 = x125 & n9557;
  assign n20297 = ~n20295 & ~n20296;
  assign n20298 = x124 & n9005;
  assign n20299 = n20297 & ~n20298;
  assign n20300 = ~n20294 & n20299;
  assign n20301 = n20300 ^ x59;
  assign n20291 = n20231 ^ n20214;
  assign n20292 = ~n20232 & n20291;
  assign n20293 = n20292 ^ n20214;
  assign n20302 = n20301 ^ n20293;
  assign n20282 = n9387 & n9878;
  assign n20283 = x120 & n9888;
  assign n20284 = x121 & n9881;
  assign n20285 = ~n20283 & ~n20284;
  assign n20286 = x122 & n10501;
  assign n20287 = n20285 & ~n20286;
  assign n20288 = ~n20282 & n20287;
  assign n20289 = n20288 ^ x62;
  assign n20274 = n7964 ^ x119;
  assign n20275 = x119 ^ x63;
  assign n20276 = n20275 ^ x119;
  assign n20277 = n20274 & n20276;
  assign n20278 = n20277 ^ x119;
  assign n20279 = ~n10177 & n20278;
  assign n20280 = n20279 ^ x119;
  assign n20266 = x117 ^ x53;
  assign n20267 = x118 ^ x116;
  assign n20268 = ~n12123 & n20267;
  assign n20269 = n20268 ^ x116;
  assign n20270 = n20269 ^ x117;
  assign n20271 = ~n20266 & n20270;
  assign n20272 = n20271 ^ x117;
  assign n20273 = ~n12893 & n20272;
  assign n20281 = n20280 ^ n20273;
  assign n20290 = n20289 ^ n20281;
  assign n20303 = n20302 ^ n20290;
  assign n20263 = n20244 ^ n20233;
  assign n20264 = n20245 & ~n20263;
  assign n20265 = n20264 ^ n20236;
  assign n20304 = n20303 ^ n20265;
  assign n20257 = n8171 & ~n10281;
  assign n20258 = x126 & n8181;
  assign n20259 = x127 & n8174;
  assign n20260 = ~n20258 & ~n20259;
  assign n20261 = ~n20257 & n20260;
  assign n20262 = n20261 ^ x56;
  assign n20305 = n20304 ^ n20262;
  assign n20322 = n20321 ^ n20305;
  assign n20380 = ~n20305 & ~n20308;
  assign n20381 = ~n20309 & ~n20380;
  assign n20382 = ~n20307 & n20381;
  assign n20383 = ~n20305 & ~n20306;
  assign n20384 = ~n20311 & ~n20383;
  assign n20385 = ~n20204 & n20384;
  assign n20386 = n20305 & n20312;
  assign n20387 = ~n20385 & ~n20386;
  assign n20388 = ~n20382 & n20387;
  assign n20369 = n9002 & ~n10570;
  assign n20370 = x124 & n9012;
  assign n20371 = x125 & n9005;
  assign n20372 = ~n20370 & ~n20371;
  assign n20373 = x126 & n9557;
  assign n20374 = n20372 & ~n20373;
  assign n20375 = ~n20369 & n20374;
  assign n20376 = n20375 ^ x59;
  assign n20359 = n9691 & n9878;
  assign n20360 = x121 & n9888;
  assign n20361 = x123 & n10501;
  assign n20362 = ~n20360 & ~n20361;
  assign n20363 = x122 & n9881;
  assign n20364 = n20362 & ~n20363;
  assign n20365 = ~n20359 & n20364;
  assign n20366 = n20365 ^ x62;
  assign n20337 = n10177 ^ x119;
  assign n20338 = x120 ^ x119;
  assign n20339 = n20338 ^ x120;
  assign n20340 = n20339 ^ n20337;
  assign n20341 = x118 ^ x63;
  assign n20342 = x118 & n20341;
  assign n20343 = n20342 ^ x120;
  assign n20344 = n20343 ^ x118;
  assign n20345 = n20340 & ~n20344;
  assign n20346 = n20345 ^ n20342;
  assign n20347 = n20346 ^ x118;
  assign n20348 = ~n20337 & n20347;
  assign n20349 = ~x118 & x119;
  assign n20350 = n20349 ^ n8244;
  assign n20351 = n20350 ^ n8244;
  assign n20352 = n8244 ^ x63;
  assign n20353 = n20352 ^ n8244;
  assign n20354 = n20351 & n20353;
  assign n20355 = n20354 ^ n8244;
  assign n20356 = ~n10177 & n20355;
  assign n20357 = n20356 ^ n8244;
  assign n20358 = ~n20348 & ~n20357;
  assign n20367 = n20366 ^ n20358;
  assign n20334 = n20289 ^ n20273;
  assign n20335 = n20281 & ~n20334;
  assign n20336 = n20335 ^ n20289;
  assign n20368 = n20367 ^ n20336;
  assign n20377 = n20376 ^ n20368;
  assign n20331 = n20303 ^ n20262;
  assign n20332 = ~n20304 & n20331;
  assign n20333 = n20332 ^ n20265;
  assign n20378 = n20377 ^ n20333;
  assign n20326 = n8171 & n11409;
  assign n20327 = x127 & n8181;
  assign n20328 = ~n20326 & ~n20327;
  assign n20329 = n20328 ^ x56;
  assign n20323 = n20301 ^ n20290;
  assign n20324 = n20302 & n20323;
  assign n20325 = n20324 ^ n20293;
  assign n20330 = n20329 ^ n20325;
  assign n20379 = n20378 ^ n20330;
  assign n20389 = n20388 ^ n20379;
  assign n20425 = ~n20325 & ~n20329;
  assign n20426 = n20388 & ~n20425;
  assign n20427 = n20325 & n20329;
  assign n20428 = n20427 ^ n20377;
  assign n20429 = n20378 & ~n20428;
  assign n20430 = n20429 ^ n20333;
  assign n20431 = n20426 & n20430;
  assign n20432 = n20425 ^ n20333;
  assign n20433 = n20377 ^ n20329;
  assign n20434 = n20433 ^ n20325;
  assign n20435 = n20427 & n20434;
  assign n20436 = n20435 ^ n20434;
  assign n20437 = ~n20432 & ~n20436;
  assign n20438 = n20437 ^ n20333;
  assign n20439 = ~n20388 & ~n20438;
  assign n20440 = n20427 ^ n20425;
  assign n20441 = n20377 & n20440;
  assign n20442 = n20441 ^ n20425;
  assign n20443 = ~n20378 & n20442;
  assign n20444 = ~n20439 & ~n20443;
  assign n20445 = ~n20431 & n20444;
  assign n20415 = n9002 & ~n10855;
  assign n20416 = x125 & n9012;
  assign n20417 = x127 & n9557;
  assign n20418 = ~n20416 & ~n20417;
  assign n20419 = x126 & n9005;
  assign n20420 = n20418 & ~n20419;
  assign n20421 = ~n20415 & n20420;
  assign n20422 = n20421 ^ x59;
  assign n20412 = n20376 ^ n20336;
  assign n20413 = ~n20368 & n20412;
  assign n20414 = n20413 ^ n20376;
  assign n20423 = n20422 ^ n20414;
  assign n20402 = n9878 & n9999;
  assign n20403 = x122 & n9888;
  assign n20404 = x123 & n9881;
  assign n20405 = ~n20403 & ~n20404;
  assign n20406 = x124 & n10501;
  assign n20407 = n20405 & ~n20406;
  assign n20408 = ~n20402 & n20407;
  assign n20409 = n20408 ^ x62;
  assign n20392 = x121 ^ x63;
  assign n20393 = n20392 ^ x121;
  assign n20394 = x121 ^ x120;
  assign n20395 = n20394 ^ x121;
  assign n20396 = n20393 & n20395;
  assign n20397 = n20396 ^ x121;
  assign n20398 = ~n10177 & n20397;
  assign n20399 = n20398 ^ x121;
  assign n20400 = n20399 ^ x56;
  assign n20401 = n20400 ^ n20280;
  assign n20410 = n20409 ^ n20401;
  assign n20390 = n20358 & ~n20366;
  assign n20391 = n20390 ^ n20357;
  assign n20411 = n20410 ^ n20391;
  assign n20424 = n20423 ^ n20411;
  assign n20446 = n20445 ^ n20424;
  assign n20479 = ~n20333 & ~n20377;
  assign n20480 = ~n20424 & ~n20479;
  assign n20481 = ~n20427 & ~n20480;
  assign n20482 = ~n20426 & n20481;
  assign n20483 = n20333 & n20377;
  assign n20484 = ~n20424 & ~n20425;
  assign n20485 = ~n20483 & ~n20484;
  assign n20486 = ~n20388 & n20485;
  assign n20487 = n20424 & ~n20430;
  assign n20488 = ~n20486 & ~n20487;
  assign n20489 = ~n20482 & n20488;
  assign n20471 = n9002 & ~n10281;
  assign n20472 = x127 & n9005;
  assign n20473 = x126 & n9012;
  assign n20474 = ~n20472 & ~n20473;
  assign n20475 = ~n20471 & n20474;
  assign n20476 = n20475 ^ x59;
  assign n20460 = n9878 & n10303;
  assign n20461 = x123 & n9888;
  assign n20462 = x124 & n9881;
  assign n20463 = ~n20461 & ~n20462;
  assign n20464 = x125 & n10501;
  assign n20465 = n20463 & ~n20464;
  assign n20466 = ~n20460 & n20465;
  assign n20467 = n20466 ^ x62;
  assign n20456 = n20280 ^ x56;
  assign n20457 = n20399 ^ n20280;
  assign n20458 = ~n20456 & ~n20457;
  assign n20459 = n20458 ^ x56;
  assign n20468 = n20467 ^ n20459;
  assign n20453 = x122 & n10177;
  assign n20454 = x121 & n12123;
  assign n20455 = ~n20453 & ~n20454;
  assign n20469 = n20468 ^ n20455;
  assign n20450 = n20409 ^ n20391;
  assign n20451 = ~n20410 & ~n20450;
  assign n20452 = n20451 ^ n20391;
  assign n20470 = n20469 ^ n20452;
  assign n20477 = n20476 ^ n20470;
  assign n20447 = n20422 ^ n20411;
  assign n20448 = n20423 & n20447;
  assign n20449 = n20448 ^ n20414;
  assign n20478 = n20477 ^ n20449;
  assign n20490 = n20489 ^ n20478;
  assign n20529 = n9002 & n11409;
  assign n20530 = x127 & n9012;
  assign n20531 = ~n20529 & ~n20530;
  assign n20532 = n20531 ^ x59;
  assign n20526 = n20476 ^ n20452;
  assign n20527 = ~n20470 & ~n20526;
  assign n20528 = n20527 ^ n20476;
  assign n20533 = n20532 ^ n20528;
  assign n20505 = n20454 ^ x123;
  assign n20506 = n20505 ^ n20454;
  assign n20507 = n20454 ^ n10177;
  assign n20508 = n20507 ^ n20454;
  assign n20509 = ~n20506 & n20508;
  assign n20510 = n20509 ^ n20454;
  assign n20511 = x122 & n20510;
  assign n20512 = n20511 ^ n20454;
  assign n20513 = n10177 ^ x122;
  assign n20514 = n9080 ^ x123;
  assign n20515 = n20514 ^ n20513;
  assign n20516 = ~x121 & ~n20392;
  assign n20517 = n20516 ^ x123;
  assign n20518 = n20517 ^ x121;
  assign n20519 = n20515 & ~n20518;
  assign n20520 = n20519 ^ n20516;
  assign n20521 = n20520 ^ x121;
  assign n20522 = n20513 & ~n20521;
  assign n20523 = ~n20512 & ~n20522;
  assign n20502 = n20459 ^ n20455;
  assign n20503 = n20468 & n20502;
  assign n20504 = n20503 ^ n20467;
  assign n20524 = n20523 ^ n20504;
  assign n20494 = n9878 & ~n10570;
  assign n20495 = x124 & n9888;
  assign n20496 = x125 & n9881;
  assign n20497 = ~n20495 & ~n20496;
  assign n20498 = x126 & n10501;
  assign n20499 = n20497 & ~n20498;
  assign n20500 = ~n20494 & n20499;
  assign n20501 = n20500 ^ x62;
  assign n20525 = n20524 ^ n20501;
  assign n20534 = n20533 ^ n20525;
  assign n20491 = n20489 ^ n20449;
  assign n20492 = ~n20478 & n20491;
  assign n20493 = n20492 ^ n20489;
  assign n20535 = n20534 ^ n20493;
  assign n20558 = n20528 & n20532;
  assign n20559 = ~n20501 & ~n20524;
  assign n20560 = n20558 & ~n20559;
  assign n20561 = ~n20528 & ~n20532;
  assign n20562 = n20501 & n20524;
  assign n20563 = n20561 & ~n20562;
  assign n20564 = ~n20560 & ~n20563;
  assign n20565 = ~n20525 & ~n20564;
  assign n20568 = ~n20561 & n20562;
  assign n20569 = ~n20560 & ~n20568;
  assign n20566 = ~n20558 & n20559;
  assign n20567 = ~n20563 & ~n20566;
  assign n20570 = n20569 ^ n20567;
  assign n20571 = ~n20493 & n20570;
  assign n20572 = n20571 ^ n20569;
  assign n20573 = ~n20565 & n20572;
  assign n20548 = n9878 & ~n10855;
  assign n20549 = x125 & n9888;
  assign n20550 = x127 & n10501;
  assign n20551 = ~n20549 & ~n20550;
  assign n20552 = x126 & n9881;
  assign n20553 = n20551 & ~n20552;
  assign n20554 = ~n20548 & n20553;
  assign n20555 = n20554 ^ x62;
  assign n20538 = x124 ^ x123;
  assign n20539 = n20538 ^ x63;
  assign n20540 = n20539 ^ n20538;
  assign n20541 = n20538 ^ n9080;
  assign n20542 = n20541 ^ n20538;
  assign n20543 = n20540 & n20542;
  assign n20544 = n20543 ^ n20538;
  assign n20545 = ~n10177 & n20544;
  assign n20546 = n20545 ^ n20538;
  assign n20547 = n20546 ^ x59;
  assign n20556 = n20555 ^ n20547;
  assign n20536 = n20504 & n20523;
  assign n20537 = n20536 ^ n20522;
  assign n20557 = n20556 ^ n20537;
  assign n20574 = n20573 ^ n20557;
  assign n20598 = n20557 & ~n20561;
  assign n20599 = ~n20562 & ~n20598;
  assign n20600 = ~n20557 & ~n20558;
  assign n20601 = ~n20566 & ~n20600;
  assign n20602 = ~n20599 & n20601;
  assign n20603 = ~n20493 & ~n20602;
  assign n20604 = n20559 & ~n20598;
  assign n20605 = ~n20568 & n20600;
  assign n20606 = ~n20604 & ~n20605;
  assign n20607 = ~n20603 & n20606;
  assign n20589 = n9878 & ~n10281;
  assign n20590 = x127 & n9881;
  assign n20591 = x126 & n9888;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = ~n20589 & n20592;
  assign n20594 = n20593 ^ x62;
  assign n20581 = x123 ^ x59;
  assign n20582 = x124 ^ x122;
  assign n20583 = ~n12123 & n20582;
  assign n20584 = n20583 ^ x122;
  assign n20585 = n20584 ^ x123;
  assign n20586 = ~n20581 & n20585;
  assign n20587 = n20586 ^ x123;
  assign n20588 = ~n12893 & n20587;
  assign n20595 = n20594 ^ n20588;
  assign n20578 = x124 & n12123;
  assign n20579 = x125 & n10177;
  assign n20580 = ~n20578 & ~n20579;
  assign n20596 = n20595 ^ n20580;
  assign n20575 = n20555 ^ n20537;
  assign n20576 = ~n20556 & n20575;
  assign n20577 = n20576 ^ n20537;
  assign n20597 = n20596 ^ n20577;
  assign n20608 = n20607 ^ n20597;
  assign n20622 = n9878 & n11409;
  assign n20623 = x127 & n9888;
  assign n20624 = ~n20622 & ~n20623;
  assign n20615 = n10302 & n12123;
  assign n20616 = x126 ^ x125;
  assign n20617 = n20616 ^ x63;
  assign n20618 = n20617 ^ x63;
  assign n20619 = n10177 & ~n20618;
  assign n20620 = n20619 ^ x63;
  assign n20621 = ~n20615 & n20620;
  assign n20625 = n20624 ^ n20621;
  assign n20612 = n20588 ^ n20580;
  assign n20613 = ~n20595 & ~n20612;
  assign n20614 = n20613 ^ n20594;
  assign n20626 = n20625 ^ n20614;
  assign n20609 = n20607 ^ n20596;
  assign n20610 = n20597 & ~n20609;
  assign n20611 = n20610 ^ n20577;
  assign n20627 = n20626 ^ n20611;
  assign n20650 = n20624 ^ x125;
  assign n20651 = ~n10302 & n20650;
  assign n20652 = n20651 ^ x125;
  assign n20653 = n20652 ^ x63;
  assign n20654 = n20653 ^ n20652;
  assign n20646 = n20624 ^ x126;
  assign n20655 = ~n20616 & n20646;
  assign n20656 = n20655 ^ x126;
  assign n20657 = n20656 ^ n20652;
  assign n20658 = ~n20654 & n20657;
  assign n20659 = n20658 ^ n20652;
  assign n20647 = n20616 & ~n20646;
  assign n20648 = x63 & n20647;
  assign n20649 = n20648 ^ n20624;
  assign n20660 = n20659 ^ n20649;
  assign n20661 = x62 & ~n20660;
  assign n20662 = n20661 ^ n20649;
  assign n20631 = x127 ^ x125;
  assign n20632 = n20631 ^ x63;
  assign n20633 = n20632 ^ x63;
  assign n20634 = n20633 ^ x62;
  assign n20635 = n20634 ^ x63;
  assign n20636 = n20635 ^ n20633;
  assign n20637 = n20633 ^ x63;
  assign n20638 = n20637 ^ n20633;
  assign n20639 = x126 ^ x124;
  assign n20640 = n20639 ^ n20633;
  assign n20641 = n20640 ^ n20633;
  assign n20642 = n20638 & n20641;
  assign n20643 = n20642 ^ n20633;
  assign n20644 = ~n20636 & n20643;
  assign n20645 = n20644 ^ n20634;
  assign n20663 = n20662 ^ n20645;
  assign n20628 = n20614 ^ n20611;
  assign n20629 = n20626 & n20628;
  assign n20630 = n20629 ^ n20611;
  assign n20664 = n20663 ^ n20630;
  assign n20668 = x127 ^ x62;
  assign n20669 = n20631 ^ x125;
  assign n20670 = x124 & x126;
  assign n20671 = n20670 ^ x125;
  assign n20672 = n20669 & n20671;
  assign n20673 = n20672 ^ x125;
  assign n20674 = ~n20668 & ~n20673;
  assign n20675 = n20674 ^ x62;
  assign n20676 = x63 & ~n20675;
  assign n20677 = n10279 & n20578;
  assign n20678 = x125 & x127;
  assign n20679 = n14116 & n20678;
  assign n20680 = ~n20677 & ~n20679;
  assign n20681 = ~n20676 & n20680;
  assign n20665 = n20662 ^ n20630;
  assign n20666 = ~n20663 & n20665;
  assign n20667 = n20666 ^ n20630;
  assign n20682 = n20681 ^ n20667;
  assign y0 = n129;
  assign y1 = n132;
  assign y2 = n148;
  assign y3 = n176;
  assign y4 = n206;
  assign y5 = ~n258;
  assign y6 = ~n303;
  assign y7 = n371;
  assign y8 = ~n432;
  assign y9 = ~n491;
  assign y10 = ~n549;
  assign y11 = ~n629;
  assign y12 = n697;
  assign y13 = ~n765;
  assign y14 = ~n847;
  assign y15 = ~n928;
  assign y16 = ~n1014;
  assign y17 = ~n1126;
  assign y18 = n1219;
  assign y19 = n1313;
  assign y20 = n1434;
  assign y21 = ~n1537;
  assign y22 = ~n1644;
  assign y23 = ~n1778;
  assign y24 = n1897;
  assign y25 = n2017;
  assign y26 = ~n2154;
  assign y27 = ~n2283;
  assign y28 = ~n2421;
  assign y29 = ~n2581;
  assign y30 = n2728;
  assign y31 = n2878;
  assign y32 = n3047;
  assign y33 = ~n3213;
  assign y34 = ~n3383;
  assign y35 = ~n3562;
  assign y36 = n3733;
  assign y37 = n3912;
  assign y38 = n4115;
  assign y39 = ~n4302;
  assign y40 = ~n4485;
  assign y41 = n4694;
  assign y42 = n4888;
  assign y43 = n5089;
  assign y44 = n5319;
  assign y45 = ~n5538;
  assign y46 = ~n5766;
  assign y47 = ~n6002;
  assign y48 = n6226;
  assign y49 = n6452;
  assign y50 = n6705;
  assign y51 = ~n6945;
  assign y52 = n7192;
  assign y53 = ~n7457;
  assign y54 = n7707;
  assign y55 = n7959;
  assign y56 = ~n8232;
  assign y57 = ~n8516;
  assign y58 = ~n8782;
  assign y59 = n9077;
  assign y60 = n9356;
  assign y61 = n9650;
  assign y62 = n9962;
  assign y63 = ~n10264;
  assign y64 = n10560;
  assign y65 = ~n10848;
  assign y66 = ~n11120;
  assign y67 = ~n11396;
  assign y68 = n11681;
  assign y69 = ~n11959;
  assign y70 = ~n12224;
  assign y71 = n12488;
  assign y72 = ~n12771;
  assign y73 = ~n13027;
  assign y74 = n13281;
  assign y75 = n13521;
  assign y76 = n13756;
  assign y77 = ~n13997;
  assign y78 = ~n14249;
  assign y79 = ~n14481;
  assign y80 = n14730;
  assign y81 = ~n14968;
  assign y82 = ~n15192;
  assign y83 = ~n15428;
  assign y84 = n15637;
  assign y85 = ~n15842;
  assign y86 = n16042;
  assign y87 = ~n16235;
  assign y88 = ~n16423;
  assign y89 = ~n16629;
  assign y90 = n16815;
  assign y91 = n16995;
  assign y92 = ~n17182;
  assign y93 = n17341;
  assign y94 = ~n17510;
  assign y95 = ~n17686;
  assign y96 = n17851;
  assign y97 = n17995;
  assign y98 = ~n18156;
  assign y99 = n18315;
  assign y100 = n18445;
  assign y101 = n18591;
  assign y102 = ~n18712;
  assign y103 = n18850;
  assign y104 = n18971;
  assign y105 = ~n19093;
  assign y106 = ~n19200;
  assign y107 = ~n19311;
  assign y108 = n19444;
  assign y109 = n19539;
  assign y110 = ~n19653;
  assign y111 = n19761;
  assign y112 = n19859;
  assign y113 = n19950;
  assign y114 = n20051;
  assign y115 = n20119;
  assign y116 = n20201;
  assign y117 = n20256;
  assign y118 = n20322;
  assign y119 = ~n20389;
  assign y120 = n20446;
  assign y121 = ~n20490;
  assign y122 = ~n20535;
  assign y123 = ~n20574;
  assign y124 = ~n20608;
  assign y125 = n20627;
  assign y126 = ~n20664;
  assign y127 = ~n20682;
endmodule