module my_module();
    logic [4:0] my_constant = 5'b11001;  // Vettore di bit di costante

    logic [4:0] my_signal;
    assign my_signal = my_constant;
  
endmodule
