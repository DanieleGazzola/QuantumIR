module Xor(input logic a, b,
           output logic xor);

    assign xor = a ^ b;
    
endmodule