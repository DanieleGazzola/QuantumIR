module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012;
  assign n129 = ~x124 & ~x125;
  assign n130 = ~x126 & n129;
  assign n131 = x126 & ~x127;
  assign n132 = ~n130 & ~n131;
  assign n133 = ~x126 & ~x127;
  assign n134 = ~x122 & ~x123;
  assign n135 = x124 & ~n134;
  assign n136 = x124 & ~x125;
  assign n137 = n131 & n136;
  assign n138 = ~n135 & ~n137;
  assign n139 = ~x124 & n134;
  assign n140 = ~x125 & x126;
  assign n141 = x127 & ~n140;
  assign n142 = n139 & ~n141;
  assign n143 = x126 ^ x125;
  assign n144 = x127 & n143;
  assign n145 = n144 ^ x125;
  assign n146 = ~n130 & ~n145;
  assign n147 = ~n142 & ~n146;
  assign n148 = x122 & ~x123;
  assign n149 = n147 & n148;
  assign n150 = ~x120 & ~x121;
  assign n151 = ~x122 & n150;
  assign n152 = n151 ^ n132;
  assign n153 = n147 ^ x123;
  assign n154 = n153 ^ n132;
  assign n155 = n152 & ~n154;
  assign n156 = n155 ^ n132;
  assign n157 = ~n149 & ~n156;
  assign n158 = ~x126 & ~n136;
  assign n159 = n158 ^ x126;
  assign n160 = n157 & n159;
  assign n161 = n160 ^ x126;
  assign n162 = ~n138 & n161;
  assign n163 = ~x125 & n157;
  assign n164 = n134 ^ x126;
  assign n165 = ~x124 & ~n164;
  assign n166 = ~x125 & ~n165;
  assign n167 = x127 & ~n166;
  assign n168 = n163 & n167;
  assign n172 = x125 & ~x126;
  assign n173 = ~n134 & ~n172;
  assign n174 = ~x124 & x127;
  assign n175 = ~n173 & n174;
  assign n169 = x125 & n134;
  assign n170 = x127 ^ x124;
  assign n171 = n169 & ~n170;
  assign n176 = n175 ^ n171;
  assign n177 = ~n157 & n176;
  assign n178 = n177 ^ n171;
  assign n179 = ~n168 & ~n178;
  assign n180 = ~n162 & n179;
  assign n192 = ~n139 & ~n163;
  assign n193 = ~x127 & ~n129;
  assign n194 = ~n192 & n193;
  assign n195 = x126 & ~n157;
  assign n196 = x125 & n135;
  assign n197 = ~n195 & n196;
  assign n198 = ~n194 & ~n197;
  assign n199 = n167 ^ n157;
  assign n200 = x126 & ~n134;
  assign n201 = ~x124 & ~n200;
  assign n202 = x125 & n201;
  assign n203 = n202 ^ n167;
  assign n204 = n203 ^ n202;
  assign n205 = n202 ^ n158;
  assign n206 = ~n204 & n205;
  assign n207 = n206 ^ n202;
  assign n208 = n199 & ~n207;
  assign n209 = n208 ^ n157;
  assign n210 = n198 & ~n209;
  assign n221 = x120 & ~x121;
  assign n222 = ~n210 & n221;
  assign n224 = ~x118 & ~x119;
  assign n225 = ~x120 & n224;
  assign n223 = n210 ^ x121;
  assign n226 = n225 ^ n223;
  assign n227 = n223 ^ n147;
  assign n228 = n226 & n227;
  assign n229 = n228 ^ n223;
  assign n230 = ~n222 & ~n229;
  assign n231 = n230 ^ n132;
  assign n232 = n150 ^ n147;
  assign n233 = ~n210 & n232;
  assign n234 = n233 ^ n147;
  assign n235 = n234 ^ x122;
  assign n236 = n235 ^ n230;
  assign n237 = ~n231 & ~n236;
  assign n238 = n237 ^ n132;
  assign n182 = n147 ^ n132;
  assign n183 = n182 ^ n147;
  assign n184 = n183 ^ n182;
  assign n185 = n182 ^ n150;
  assign n186 = ~n184 & n185;
  assign n187 = n186 ^ n182;
  assign n188 = ~x122 & n187;
  assign n189 = n188 ^ n182;
  assign n181 = ~x122 & n147;
  assign n190 = n189 ^ n181;
  assign n191 = n189 ^ n152;
  assign n211 = n210 ^ n189;
  assign n212 = ~n189 & n211;
  assign n213 = n212 ^ n189;
  assign n214 = n191 & ~n213;
  assign n215 = n214 ^ n212;
  assign n216 = n215 ^ n189;
  assign n217 = n216 ^ n210;
  assign n218 = n190 & n217;
  assign n219 = n218 ^ n181;
  assign n220 = n219 ^ x123;
  assign n239 = n238 ^ n220;
  assign n240 = n220 ^ n133;
  assign n241 = ~n239 & n240;
  assign n242 = n241 ^ n220;
  assign n243 = n180 & ~n242;
  assign n252 = x118 & ~x119;
  assign n253 = ~n243 & n252;
  assign n254 = n243 ^ x119;
  assign n255 = n254 ^ n210;
  assign n256 = ~x116 & ~x117;
  assign n257 = ~x118 & n256;
  assign n258 = n257 ^ n254;
  assign n259 = ~n255 & n258;
  assign n260 = n259 ^ n254;
  assign n261 = ~n253 & ~n260;
  assign n262 = n261 ^ n147;
  assign n263 = n224 ^ n210;
  assign n264 = ~n243 & ~n263;
  assign n265 = n264 ^ n210;
  assign n266 = n265 ^ x120;
  assign n267 = n266 ^ n261;
  assign n268 = ~n262 & n267;
  assign n269 = n268 ^ n147;
  assign n270 = n269 ^ n132;
  assign n279 = ~x120 & ~n210;
  assign n271 = n210 ^ n147;
  assign n272 = n271 ^ n210;
  assign n273 = n272 ^ n271;
  assign n274 = n271 ^ n224;
  assign n275 = n273 & ~n274;
  assign n276 = n275 ^ n271;
  assign n277 = ~x120 & ~n276;
  assign n278 = n277 ^ n271;
  assign n280 = n279 ^ n278;
  assign n281 = n225 ^ n224;
  assign n282 = ~n147 & ~n281;
  assign n283 = n282 ^ n224;
  assign n284 = n283 ^ n278;
  assign n285 = n278 ^ n243;
  assign n286 = n278 & ~n285;
  assign n287 = n286 ^ n278;
  assign n288 = n284 & n287;
  assign n289 = n288 ^ n286;
  assign n290 = n289 ^ n278;
  assign n291 = n290 ^ n243;
  assign n292 = ~n280 & ~n291;
  assign n293 = n292 ^ n279;
  assign n294 = n293 ^ x121;
  assign n295 = n294 ^ n269;
  assign n296 = n270 & n295;
  assign n297 = n296 ^ n132;
  assign n247 = ~n231 & ~n243;
  assign n248 = n247 ^ n235;
  assign n348 = ~n133 & n248;
  assign n244 = n220 ^ n180;
  assign n245 = ~n238 & ~n244;
  assign n246 = n245 ^ n220;
  assign n249 = n248 ^ n246;
  assign n250 = ~n133 & n249;
  assign n251 = n250 ^ n248;
  assign n349 = n348 ^ n251;
  assign n350 = n297 & n349;
  assign n351 = n350 ^ n251;
  assign n298 = ~n133 & ~n248;
  assign n299 = ~n297 & ~n298;
  assign n300 = ~n251 & ~n299;
  assign n301 = n256 ^ n243;
  assign n302 = ~n300 & ~n301;
  assign n303 = n302 ^ n243;
  assign n304 = n303 ^ x118;
  assign n305 = n304 ^ n210;
  assign n306 = x116 & ~x117;
  assign n307 = ~n300 & n306;
  assign n308 = n300 ^ x117;
  assign n309 = n308 ^ n243;
  assign n310 = ~x114 & ~x115;
  assign n311 = ~x116 & n310;
  assign n312 = n311 ^ n308;
  assign n313 = ~n309 & n312;
  assign n314 = n313 ^ n308;
  assign n315 = ~n307 & ~n314;
  assign n316 = n315 ^ n304;
  assign n317 = ~n305 & n316;
  assign n318 = n317 ^ n210;
  assign n319 = n318 ^ n147;
  assign n328 = ~x118 & ~n243;
  assign n320 = n243 ^ n210;
  assign n321 = n320 ^ n243;
  assign n322 = n321 ^ n320;
  assign n323 = n320 ^ n256;
  assign n324 = n322 & n323;
  assign n325 = n324 ^ n320;
  assign n326 = ~x118 & n325;
  assign n327 = n326 ^ n320;
  assign n329 = n328 ^ n327;
  assign n330 = n257 ^ n256;
  assign n331 = n210 & ~n330;
  assign n332 = n331 ^ n256;
  assign n333 = n332 ^ n327;
  assign n334 = n327 ^ n300;
  assign n335 = ~n327 & n334;
  assign n336 = n335 ^ n327;
  assign n337 = ~n333 & ~n336;
  assign n338 = n337 ^ n335;
  assign n339 = n338 ^ n327;
  assign n340 = n339 ^ n300;
  assign n341 = n329 & n340;
  assign n342 = n341 ^ n328;
  assign n343 = n342 ^ x119;
  assign n344 = n343 ^ n318;
  assign n345 = ~n319 & ~n344;
  assign n346 = n345 ^ n147;
  assign n347 = n346 ^ n132;
  assign n354 = ~n262 & ~n300;
  assign n355 = n354 ^ n266;
  assign n356 = n355 ^ n346;
  assign n357 = n347 & ~n356;
  assign n358 = n357 ^ n132;
  assign n352 = n270 & ~n300;
  assign n353 = n352 ^ n294;
  assign n359 = n358 ^ n353;
  assign n360 = n353 ^ n133;
  assign n361 = ~n359 & n360;
  assign n362 = n361 ^ n353;
  assign n363 = ~n351 & ~n362;
  assign n366 = n310 ^ n300;
  assign n367 = ~n363 & ~n366;
  assign n368 = n367 ^ n300;
  assign n369 = n368 ^ x116;
  assign n370 = n369 ^ n243;
  assign n371 = x114 & ~x115;
  assign n372 = ~n363 & n371;
  assign n373 = n363 ^ x115;
  assign n374 = n373 ^ n300;
  assign n375 = ~x112 & ~x113;
  assign n376 = ~x114 & n375;
  assign n377 = n376 ^ n373;
  assign n378 = ~n374 & n377;
  assign n379 = n378 ^ n373;
  assign n380 = ~n372 & ~n379;
  assign n381 = n380 ^ n369;
  assign n382 = ~n370 & n381;
  assign n383 = n382 ^ n243;
  assign n384 = n383 ^ n210;
  assign n393 = ~x116 & ~n300;
  assign n385 = n300 ^ n243;
  assign n386 = n385 ^ n300;
  assign n387 = n386 ^ n385;
  assign n388 = n385 ^ n310;
  assign n389 = n387 & n388;
  assign n390 = n389 ^ n385;
  assign n391 = ~x116 & n390;
  assign n392 = n391 ^ n385;
  assign n394 = n393 ^ n392;
  assign n395 = n311 ^ n310;
  assign n396 = n243 & ~n395;
  assign n397 = n396 ^ n310;
  assign n398 = n397 ^ n392;
  assign n399 = n392 ^ n363;
  assign n400 = ~n392 & n399;
  assign n401 = n400 ^ n392;
  assign n402 = ~n398 & ~n401;
  assign n403 = n402 ^ n400;
  assign n404 = n403 ^ n392;
  assign n405 = n404 ^ n363;
  assign n406 = n394 & n405;
  assign n407 = n406 ^ n393;
  assign n408 = n407 ^ x117;
  assign n409 = n408 ^ n383;
  assign n410 = n384 & ~n409;
  assign n411 = n410 ^ n210;
  assign n412 = n411 ^ n147;
  assign n413 = n315 ^ n210;
  assign n414 = ~n363 & n413;
  assign n415 = n414 ^ n304;
  assign n416 = n415 ^ n411;
  assign n417 = ~n412 & n416;
  assign n418 = n417 ^ n147;
  assign n419 = n418 ^ n132;
  assign n420 = ~n319 & ~n363;
  assign n421 = n420 ^ n343;
  assign n422 = n421 ^ n418;
  assign n423 = n419 & n422;
  assign n424 = n423 ^ n132;
  assign n364 = n347 & ~n363;
  assign n365 = n364 ^ n355;
  assign n426 = n424 ^ n365;
  assign n425 = n365 & n424;
  assign n427 = n426 ^ n425;
  assign n428 = ~n353 & n363;
  assign n429 = ~n359 & n428;
  assign n430 = n429 ^ n359;
  assign n431 = n430 ^ n425;
  assign n432 = n431 ^ n425;
  assign n433 = n427 & n432;
  assign n434 = n433 ^ n425;
  assign n435 = ~n133 & n434;
  assign n436 = n435 ^ n425;
  assign n437 = n375 ^ n363;
  assign n438 = ~n436 & ~n437;
  assign n439 = n438 ^ n363;
  assign n440 = n439 ^ x114;
  assign n441 = n440 ^ n300;
  assign n442 = x112 & ~x113;
  assign n443 = ~n436 & n442;
  assign n444 = n436 ^ x113;
  assign n445 = n444 ^ n363;
  assign n446 = ~x110 & ~x111;
  assign n447 = ~x112 & n446;
  assign n448 = n447 ^ n444;
  assign n449 = ~n445 & n448;
  assign n450 = n449 ^ n444;
  assign n451 = ~n443 & ~n450;
  assign n452 = n451 ^ n440;
  assign n453 = ~n441 & n452;
  assign n454 = n453 ^ n300;
  assign n455 = n454 ^ n243;
  assign n464 = ~x114 & ~n363;
  assign n456 = n363 ^ n300;
  assign n457 = n456 ^ n363;
  assign n458 = n457 ^ n456;
  assign n459 = n456 ^ n375;
  assign n460 = n458 & n459;
  assign n461 = n460 ^ n456;
  assign n462 = ~x114 & n461;
  assign n463 = n462 ^ n456;
  assign n465 = n464 ^ n463;
  assign n466 = n376 ^ n375;
  assign n467 = n300 & ~n466;
  assign n468 = n467 ^ n375;
  assign n469 = n468 ^ n463;
  assign n470 = n463 ^ n436;
  assign n471 = ~n463 & n470;
  assign n472 = n471 ^ n463;
  assign n473 = ~n469 & ~n472;
  assign n474 = n473 ^ n471;
  assign n475 = n474 ^ n463;
  assign n476 = n475 ^ n436;
  assign n477 = n465 & n476;
  assign n478 = n477 ^ n464;
  assign n479 = n478 ^ x115;
  assign n480 = n479 ^ n454;
  assign n481 = n455 & ~n480;
  assign n482 = n481 ^ n243;
  assign n483 = n482 ^ n210;
  assign n484 = n380 ^ n243;
  assign n485 = ~n436 & n484;
  assign n486 = n485 ^ n369;
  assign n487 = n486 ^ n482;
  assign n488 = n483 & n487;
  assign n489 = n488 ^ n210;
  assign n490 = n489 ^ n147;
  assign n491 = n384 & ~n436;
  assign n492 = n491 ^ n408;
  assign n493 = n492 ^ n489;
  assign n494 = ~n490 & ~n493;
  assign n495 = n494 ^ n147;
  assign n496 = n495 ^ n132;
  assign n497 = ~n412 & ~n436;
  assign n498 = n497 ^ n415;
  assign n499 = n498 ^ n495;
  assign n500 = n496 & ~n499;
  assign n501 = n500 ^ n132;
  assign n502 = n419 & ~n436;
  assign n503 = n502 ^ n421;
  assign n504 = ~n501 & n503;
  assign n505 = n501 & ~n503;
  assign n506 = n505 ^ n133;
  assign n507 = n506 ^ n505;
  assign n508 = n430 ^ n365;
  assign n509 = ~n424 & n508;
  assign n510 = n509 ^ n365;
  assign n511 = n510 ^ n505;
  assign n512 = ~n507 & n511;
  assign n513 = n512 ^ n505;
  assign n514 = ~n504 & n513;
  assign n517 = n446 ^ n436;
  assign n518 = ~n514 & ~n517;
  assign n519 = n518 ^ n436;
  assign n520 = n519 ^ x112;
  assign n521 = n520 ^ n363;
  assign n522 = x110 & ~x111;
  assign n523 = ~n514 & n522;
  assign n525 = ~x108 & ~x109;
  assign n526 = ~x110 & n525;
  assign n524 = n514 ^ x111;
  assign n527 = n526 ^ n524;
  assign n528 = n524 ^ n436;
  assign n529 = n527 & ~n528;
  assign n530 = n529 ^ n524;
  assign n531 = ~n523 & ~n530;
  assign n532 = n531 ^ n520;
  assign n533 = ~n521 & n532;
  assign n534 = n533 ^ n363;
  assign n535 = n534 ^ n300;
  assign n544 = ~x112 & ~n436;
  assign n536 = n436 ^ n363;
  assign n537 = n536 ^ n436;
  assign n538 = n537 ^ n536;
  assign n539 = n536 ^ n446;
  assign n540 = n538 & n539;
  assign n541 = n540 ^ n536;
  assign n542 = ~x112 & n541;
  assign n543 = n542 ^ n536;
  assign n545 = n544 ^ n543;
  assign n546 = n447 ^ n446;
  assign n547 = n363 & ~n546;
  assign n548 = n547 ^ n446;
  assign n549 = n548 ^ n543;
  assign n550 = n543 ^ n514;
  assign n551 = ~n543 & n550;
  assign n552 = n551 ^ n543;
  assign n553 = ~n549 & ~n552;
  assign n554 = n553 ^ n551;
  assign n555 = n554 ^ n543;
  assign n556 = n555 ^ n514;
  assign n557 = n545 & n556;
  assign n558 = n557 ^ n544;
  assign n559 = n558 ^ x113;
  assign n560 = n559 ^ n534;
  assign n561 = n535 & ~n560;
  assign n562 = n561 ^ n300;
  assign n563 = n562 ^ n243;
  assign n564 = n451 ^ n300;
  assign n565 = ~n514 & n564;
  assign n566 = n565 ^ n440;
  assign n567 = n566 ^ n562;
  assign n568 = n563 & n567;
  assign n569 = n568 ^ n243;
  assign n570 = n569 ^ n210;
  assign n571 = n455 & ~n514;
  assign n572 = n571 ^ n479;
  assign n573 = n572 ^ n569;
  assign n574 = n570 & ~n573;
  assign n575 = n574 ^ n210;
  assign n576 = n575 ^ n147;
  assign n577 = n483 & ~n514;
  assign n578 = n577 ^ n486;
  assign n579 = n578 ^ n575;
  assign n580 = ~n576 & n579;
  assign n581 = n580 ^ n147;
  assign n582 = n581 ^ n132;
  assign n583 = ~n490 & ~n514;
  assign n584 = n583 ^ n492;
  assign n585 = n584 ^ n581;
  assign n586 = n582 & n585;
  assign n587 = n586 ^ n132;
  assign n589 = n510 ^ n503;
  assign n590 = ~n501 & ~n589;
  assign n591 = n590 ^ n503;
  assign n689 = ~n133 & ~n591;
  assign n515 = n496 & ~n514;
  assign n516 = n515 ^ n498;
  assign n690 = n689 ^ n516;
  assign n691 = ~n587 & n690;
  assign n692 = n691 ^ n516;
  assign n693 = n692 ^ n133;
  assign n694 = n693 ^ n692;
  assign n592 = n591 ^ n516;
  assign n593 = n592 ^ n516;
  assign n594 = n593 ^ n133;
  assign n595 = n594 ^ n593;
  assign n596 = n595 ^ n516;
  assign n588 = n587 ^ n516;
  assign n597 = n596 ^ n588;
  assign n598 = n593 ^ n587;
  assign n599 = n598 ^ n516;
  assign n600 = n599 ^ n516;
  assign n601 = ~n595 & ~n600;
  assign n602 = n601 ^ n595;
  assign n603 = n599 & ~n602;
  assign n604 = n603 ^ n516;
  assign n605 = ~n597 & ~n604;
  assign n606 = n605 ^ n601;
  assign n607 = n606 ^ n516;
  assign n608 = n607 ^ n588;
  assign n609 = n525 ^ n514;
  assign n610 = ~n608 & ~n609;
  assign n611 = n610 ^ n514;
  assign n612 = n611 ^ x110;
  assign n613 = n612 ^ n436;
  assign n614 = x108 & ~x109;
  assign n615 = ~n608 & n614;
  assign n616 = ~x106 & ~x107;
  assign n617 = ~x108 & n616;
  assign n618 = n617 ^ n514;
  assign n619 = n608 ^ x109;
  assign n620 = n619 ^ n514;
  assign n621 = ~n618 & ~n620;
  assign n622 = n621 ^ n514;
  assign n623 = ~n615 & n622;
  assign n624 = n623 ^ n612;
  assign n625 = ~n613 & n624;
  assign n626 = n625 ^ n436;
  assign n627 = n626 ^ n363;
  assign n636 = ~x110 & ~n514;
  assign n628 = n514 ^ n436;
  assign n629 = n628 ^ n514;
  assign n630 = n629 ^ n628;
  assign n631 = n628 ^ n525;
  assign n632 = n630 & n631;
  assign n633 = n632 ^ n628;
  assign n634 = ~x110 & n633;
  assign n635 = n634 ^ n628;
  assign n637 = n636 ^ n635;
  assign n638 = n526 ^ n525;
  assign n639 = n436 & ~n638;
  assign n640 = n639 ^ n525;
  assign n641 = n640 ^ n635;
  assign n642 = n635 ^ n608;
  assign n643 = ~n635 & n642;
  assign n644 = n643 ^ n635;
  assign n645 = ~n641 & ~n644;
  assign n646 = n645 ^ n643;
  assign n647 = n646 ^ n635;
  assign n648 = n647 ^ n608;
  assign n649 = n637 & n648;
  assign n650 = n649 ^ n636;
  assign n651 = n650 ^ x111;
  assign n652 = n651 ^ n626;
  assign n653 = n627 & ~n652;
  assign n654 = n653 ^ n363;
  assign n655 = n654 ^ n300;
  assign n656 = n531 ^ n363;
  assign n657 = ~n608 & n656;
  assign n658 = n657 ^ n520;
  assign n659 = n658 ^ n654;
  assign n660 = n655 & n659;
  assign n661 = n660 ^ n300;
  assign n662 = n661 ^ n243;
  assign n663 = n535 & ~n608;
  assign n664 = n663 ^ n559;
  assign n665 = n664 ^ n661;
  assign n666 = n662 & ~n665;
  assign n667 = n666 ^ n243;
  assign n668 = n667 ^ n210;
  assign n669 = n563 & ~n608;
  assign n670 = n669 ^ n566;
  assign n671 = n670 ^ n667;
  assign n672 = n668 & n671;
  assign n673 = n672 ^ n210;
  assign n674 = n673 ^ n147;
  assign n675 = n570 & ~n608;
  assign n676 = n675 ^ n572;
  assign n677 = n676 ^ n673;
  assign n678 = ~n674 & ~n677;
  assign n679 = n678 ^ n147;
  assign n680 = n679 ^ n132;
  assign n683 = ~n576 & ~n608;
  assign n684 = n683 ^ n578;
  assign n685 = n684 ^ n679;
  assign n686 = n680 & ~n685;
  assign n687 = n686 ^ n132;
  assign n695 = n694 ^ n687;
  assign n681 = n582 & ~n608;
  assign n682 = n681 ^ n584;
  assign n688 = n687 ^ n682;
  assign n696 = n695 ^ n688;
  assign n697 = n692 ^ n682;
  assign n698 = n697 ^ n687;
  assign n699 = n698 ^ n687;
  assign n700 = ~n694 & ~n699;
  assign n701 = n700 ^ n694;
  assign n702 = n698 & ~n701;
  assign n703 = n702 ^ n687;
  assign n704 = n696 & ~n703;
  assign n705 = n704 ^ n700;
  assign n706 = n705 ^ n687;
  assign n707 = n706 ^ n688;
  assign n710 = n616 ^ n608;
  assign n711 = n707 & ~n710;
  assign n712 = n711 ^ n608;
  assign n713 = n712 ^ x108;
  assign n714 = n713 ^ n514;
  assign n715 = x106 & ~x107;
  assign n716 = n707 & n715;
  assign n717 = ~x104 & ~x105;
  assign n718 = ~x106 & n717;
  assign n719 = n718 ^ n608;
  assign n720 = n707 ^ x107;
  assign n721 = n720 ^ n608;
  assign n722 = ~n719 & n721;
  assign n723 = n722 ^ n608;
  assign n724 = ~n716 & n723;
  assign n725 = n724 ^ n713;
  assign n726 = ~n714 & n725;
  assign n727 = n726 ^ n514;
  assign n728 = n727 ^ n436;
  assign n788 = ~n687 & ~n697;
  assign n789 = n788 ^ n682;
  assign n790 = ~n133 & n789;
  assign n708 = n680 & n707;
  assign n709 = n708 ^ n684;
  assign n799 = n709 ^ n133;
  assign n730 = x108 & n514;
  assign n731 = n730 ^ n618;
  assign n732 = ~n608 & ~n731;
  assign n733 = n732 ^ n618;
  assign n729 = ~x108 & ~n608;
  assign n734 = n733 ^ n729;
  assign n735 = n616 ^ n514;
  assign n736 = n735 ^ n733;
  assign n737 = n733 ^ n707;
  assign n738 = n733 & n737;
  assign n739 = n738 ^ n733;
  assign n740 = n736 & n739;
  assign n741 = n740 ^ n738;
  assign n742 = n741 ^ n733;
  assign n743 = n742 ^ n707;
  assign n744 = ~n734 & n743;
  assign n745 = n744 ^ n729;
  assign n746 = n745 ^ x109;
  assign n747 = n746 ^ n727;
  assign n748 = n728 & ~n747;
  assign n749 = n748 ^ n436;
  assign n750 = n749 ^ n363;
  assign n751 = n623 ^ n436;
  assign n752 = n707 & n751;
  assign n753 = n752 ^ n612;
  assign n754 = n753 ^ n749;
  assign n755 = n750 & n754;
  assign n756 = n755 ^ n363;
  assign n757 = n756 ^ n300;
  assign n758 = n627 & n707;
  assign n759 = n758 ^ n651;
  assign n760 = n759 ^ n756;
  assign n761 = n757 & ~n760;
  assign n762 = n761 ^ n300;
  assign n763 = n762 ^ n243;
  assign n764 = n655 & n707;
  assign n765 = n764 ^ n658;
  assign n766 = n765 ^ n762;
  assign n767 = n763 & n766;
  assign n768 = n767 ^ n243;
  assign n769 = n768 ^ n210;
  assign n770 = n662 & n707;
  assign n771 = n770 ^ n664;
  assign n772 = n771 ^ n768;
  assign n773 = n769 & ~n772;
  assign n774 = n773 ^ n210;
  assign n775 = n774 ^ n147;
  assign n776 = n668 & n707;
  assign n777 = n776 ^ n670;
  assign n778 = n777 ^ n774;
  assign n779 = ~n775 & n778;
  assign n780 = n779 ^ n147;
  assign n781 = n780 ^ n132;
  assign n782 = ~n674 & n707;
  assign n783 = n782 ^ n676;
  assign n784 = n783 ^ n780;
  assign n785 = n781 & n784;
  assign n786 = n785 ^ n132;
  assign n800 = n786 ^ n709;
  assign n801 = ~n799 & n800;
  assign n802 = n801 ^ n709;
  assign n803 = ~n790 & n802;
  assign n804 = n728 & ~n803;
  assign n805 = n804 ^ n746;
  assign n806 = ~n363 & ~n805;
  assign n807 = n750 & ~n803;
  assign n808 = n807 ^ n753;
  assign n809 = ~n300 & n808;
  assign n810 = ~n806 & ~n809;
  assign n811 = n724 ^ n514;
  assign n812 = ~n803 & n811;
  assign n813 = n812 ^ n713;
  assign n814 = n813 ^ n436;
  assign n816 = x106 & n608;
  assign n817 = n816 ^ n719;
  assign n818 = n707 & ~n817;
  assign n819 = n818 ^ n719;
  assign n815 = ~x106 & n707;
  assign n820 = n819 ^ n815;
  assign n821 = n717 ^ n608;
  assign n822 = n821 ^ n819;
  assign n823 = n819 ^ n803;
  assign n824 = n819 & ~n823;
  assign n825 = n824 ^ n819;
  assign n826 = n822 & n825;
  assign n827 = n826 ^ n824;
  assign n828 = n827 ^ n819;
  assign n829 = n828 ^ n803;
  assign n830 = ~n820 & ~n829;
  assign n831 = n830 ^ n815;
  assign n832 = n831 ^ x107;
  assign n833 = n832 ^ n514;
  assign n834 = n717 ^ n707;
  assign n835 = ~n803 & n834;
  assign n836 = n835 ^ n707;
  assign n837 = n836 ^ x106;
  assign n838 = n837 ^ n608;
  assign n839 = x104 & ~x105;
  assign n840 = ~n803 & n839;
  assign n841 = ~x102 & ~x103;
  assign n842 = ~x104 & n841;
  assign n843 = n842 ^ n707;
  assign n844 = n803 ^ x105;
  assign n845 = n844 ^ n707;
  assign n846 = n843 & n845;
  assign n847 = n846 ^ n707;
  assign n848 = ~n840 & ~n847;
  assign n849 = n848 ^ n837;
  assign n850 = n838 & ~n849;
  assign n851 = n850 ^ n608;
  assign n852 = n851 ^ n832;
  assign n853 = n833 & ~n852;
  assign n854 = n853 ^ n514;
  assign n855 = n854 ^ n813;
  assign n856 = ~n814 & n855;
  assign n857 = n856 ^ n436;
  assign n858 = n810 & n857;
  assign n859 = n808 ^ n300;
  assign n860 = n363 & n805;
  assign n861 = n860 ^ n808;
  assign n862 = ~n859 & n861;
  assign n863 = n862 ^ n300;
  assign n864 = ~n858 & ~n863;
  assign n865 = n243 & ~n864;
  assign n866 = n763 & ~n803;
  assign n867 = n866 ^ n765;
  assign n868 = n865 & ~n867;
  assign n869 = n757 & ~n803;
  assign n870 = n869 ^ n759;
  assign n871 = n870 ^ n210;
  assign n872 = n870 ^ n243;
  assign n873 = n872 ^ n243;
  assign n874 = n867 ^ n243;
  assign n875 = n873 & n874;
  assign n876 = n875 ^ n243;
  assign n877 = n871 & ~n876;
  assign n878 = n877 ^ n210;
  assign n879 = ~n864 & n878;
  assign n880 = n867 ^ n210;
  assign n881 = n243 & n870;
  assign n882 = n881 ^ n867;
  assign n883 = ~n880 & n882;
  assign n884 = n883 ^ n210;
  assign n885 = ~n879 & ~n884;
  assign n886 = ~n868 & n885;
  assign n887 = n886 ^ n147;
  assign n888 = n769 & ~n803;
  assign n889 = n888 ^ n771;
  assign n890 = n889 ^ n886;
  assign n891 = n887 & n890;
  assign n892 = n891 ^ n147;
  assign n893 = n892 ^ n132;
  assign n787 = n786 ^ n133;
  assign n791 = n790 ^ n787;
  assign n792 = n791 ^ n787;
  assign n793 = n787 ^ n786;
  assign n794 = n793 ^ n787;
  assign n795 = n792 & ~n794;
  assign n796 = n795 ^ n787;
  assign n797 = n709 & n796;
  assign n798 = n797 ^ n787;
  assign n894 = ~n775 & ~n803;
  assign n895 = n894 ^ n777;
  assign n896 = n895 ^ n892;
  assign n897 = n893 & ~n896;
  assign n898 = n897 ^ n132;
  assign n899 = n898 ^ n133;
  assign n900 = n781 & ~n803;
  assign n901 = n900 ^ n783;
  assign n902 = n901 ^ n898;
  assign n903 = ~n899 & ~n902;
  assign n904 = n903 ^ n898;
  assign n905 = ~n798 & n904;
  assign n1008 = n893 & ~n905;
  assign n1009 = n1008 ^ n895;
  assign n906 = x102 & ~n905;
  assign n907 = ~x103 & n906;
  assign n908 = ~x100 & ~x101;
  assign n909 = ~x102 & n908;
  assign n910 = n909 ^ n803;
  assign n911 = n905 ^ x103;
  assign n912 = n911 ^ n803;
  assign n913 = ~n910 & ~n912;
  assign n914 = n913 ^ n803;
  assign n915 = ~n907 & n914;
  assign n916 = n915 ^ n707;
  assign n917 = n841 ^ n803;
  assign n918 = ~n905 & ~n917;
  assign n919 = n918 ^ n803;
  assign n920 = n919 ^ x104;
  assign n921 = n920 ^ n915;
  assign n922 = ~n916 & n921;
  assign n923 = n922 ^ n707;
  assign n924 = n923 ^ n608;
  assign n926 = x104 & ~n707;
  assign n927 = n926 ^ n843;
  assign n928 = ~n803 & n927;
  assign n929 = n928 ^ n843;
  assign n925 = ~x104 & ~n803;
  assign n930 = n929 ^ n925;
  assign n931 = n841 ^ n707;
  assign n932 = n931 ^ n929;
  assign n933 = n929 ^ n905;
  assign n934 = ~n929 & n933;
  assign n935 = n934 ^ n929;
  assign n936 = n932 & ~n935;
  assign n937 = n936 ^ n934;
  assign n938 = n937 ^ n929;
  assign n939 = n938 ^ n905;
  assign n940 = n930 & n939;
  assign n941 = n940 ^ n925;
  assign n942 = n941 ^ x105;
  assign n943 = n942 ^ n923;
  assign n944 = ~n924 & n943;
  assign n945 = n944 ^ n608;
  assign n946 = n945 ^ n514;
  assign n947 = n848 ^ n608;
  assign n948 = ~n905 & n947;
  assign n949 = n948 ^ n837;
  assign n950 = n949 ^ n945;
  assign n951 = n946 & ~n950;
  assign n952 = n951 ^ n514;
  assign n953 = n952 ^ n436;
  assign n954 = n851 ^ n514;
  assign n955 = ~n905 & n954;
  assign n956 = n955 ^ n832;
  assign n957 = n956 ^ n952;
  assign n958 = n953 & ~n957;
  assign n959 = n958 ^ n436;
  assign n960 = n959 ^ n363;
  assign n961 = n854 ^ n436;
  assign n962 = ~n905 & n961;
  assign n963 = n962 ^ n813;
  assign n964 = n963 ^ n959;
  assign n965 = n960 & n964;
  assign n966 = n965 ^ n363;
  assign n967 = n966 ^ n300;
  assign n968 = n857 ^ n363;
  assign n969 = ~n905 & n968;
  assign n970 = n969 ^ n805;
  assign n971 = n970 ^ n966;
  assign n972 = n967 & ~n971;
  assign n973 = n972 ^ n300;
  assign n974 = n973 ^ n243;
  assign n975 = n857 ^ n805;
  assign n976 = n968 & ~n975;
  assign n977 = n976 ^ n363;
  assign n978 = n977 ^ n300;
  assign n979 = ~n905 & n978;
  assign n980 = n979 ^ n808;
  assign n981 = n980 ^ n973;
  assign n982 = n974 & n981;
  assign n983 = n982 ^ n243;
  assign n984 = n983 ^ n210;
  assign n985 = n864 ^ n243;
  assign n986 = ~n905 & ~n985;
  assign n987 = n986 ^ n870;
  assign n988 = n987 ^ n983;
  assign n989 = n984 & ~n988;
  assign n990 = n989 ^ n210;
  assign n991 = n990 ^ n147;
  assign n992 = n870 ^ n864;
  assign n993 = ~n985 & n992;
  assign n994 = n993 ^ n243;
  assign n995 = n994 ^ n210;
  assign n996 = ~n905 & n995;
  assign n997 = n996 ^ n867;
  assign n998 = n997 ^ n990;
  assign n999 = ~n991 & n998;
  assign n1000 = n999 ^ n147;
  assign n1001 = n1000 ^ n132;
  assign n1002 = n887 & ~n905;
  assign n1003 = n1002 ^ n889;
  assign n1004 = n1003 ^ n1000;
  assign n1005 = n1001 & n1004;
  assign n1006 = n1005 ^ n132;
  assign n1007 = n1006 ^ n133;
  assign n1010 = n1009 ^ n1007;
  assign n1011 = n899 ^ n798;
  assign n1012 = n1011 ^ n899;
  assign n1013 = n899 ^ n898;
  assign n1014 = n1013 ^ n899;
  assign n1015 = n1012 & ~n1014;
  assign n1016 = n1015 ^ n899;
  assign n1017 = ~n901 & n1016;
  assign n1018 = n1017 ^ n899;
  assign n1019 = ~n1007 & ~n1018;
  assign n1020 = n1010 & n1019;
  assign n1021 = n1020 ^ n1010;
  assign n1022 = ~x98 & ~x99;
  assign n1023 = ~x100 & n1022;
  assign n1028 = n905 ^ x101;
  assign n1024 = n1009 ^ n1006;
  assign n1025 = ~n1007 & ~n1024;
  assign n1026 = n1025 ^ n133;
  assign n1027 = ~n1018 & ~n1026;
  assign n1029 = n1028 ^ n1027;
  assign n1030 = n905 ^ x102;
  assign n1031 = n1030 ^ n1027;
  assign n1032 = n1030 ^ n905;
  assign n1033 = n1032 ^ n1030;
  assign n1034 = ~n1031 & ~n1033;
  assign n1035 = n1034 ^ n1030;
  assign n1036 = n1029 & n1035;
  assign n1037 = n1036 ^ n1030;
  assign n1038 = n1023 & n1037;
  assign n1039 = x101 & ~n905;
  assign n1040 = x100 & ~x101;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = ~x102 & ~n1041;
  assign n1043 = ~n1027 & n1042;
  assign n1044 = n803 & ~n1043;
  assign n1045 = n906 & n1027;
  assign n1046 = ~x101 & n1045;
  assign n1047 = n1044 & ~n1046;
  assign n1048 = ~n1038 & n1047;
  assign n1059 = n1027 ^ x101;
  assign n1060 = n1027 ^ n1023;
  assign n1061 = n1059 & ~n1060;
  assign n1062 = n1061 ^ n1027;
  assign n1049 = ~n905 & n1023;
  assign n1050 = n908 & ~n1049;
  assign n1051 = n1050 ^ n1023;
  assign n1052 = n1051 ^ n1050;
  assign n1053 = n1050 ^ n1039;
  assign n1054 = n1053 ^ n1050;
  assign n1055 = ~n1052 & n1054;
  assign n1056 = n1055 ^ n1050;
  assign n1057 = n1027 & n1056;
  assign n1058 = n1057 ^ n1050;
  assign n1063 = n1062 ^ n1058;
  assign n1064 = n1063 ^ n1058;
  assign n1065 = n1058 ^ n905;
  assign n1066 = n1065 ^ n1058;
  assign n1067 = n1064 & n1066;
  assign n1068 = n1067 ^ n1058;
  assign n1069 = x102 & n1068;
  assign n1070 = n1069 ^ n1058;
  assign n1071 = ~n1048 & ~n1070;
  assign n1072 = n1071 ^ n707;
  assign n1081 = ~x102 & ~n905;
  assign n1073 = n905 ^ n803;
  assign n1074 = n1073 ^ n905;
  assign n1075 = n1074 ^ n1073;
  assign n1076 = n1073 ^ n908;
  assign n1077 = n1075 & n1076;
  assign n1078 = n1077 ^ n1073;
  assign n1079 = ~x102 & n1078;
  assign n1080 = n1079 ^ n1073;
  assign n1082 = n1081 ^ n1080;
  assign n1083 = n908 ^ n803;
  assign n1084 = n1083 ^ n1080;
  assign n1085 = n1080 ^ n1027;
  assign n1086 = ~n1080 & n1085;
  assign n1087 = n1086 ^ n1080;
  assign n1088 = ~n1084 & ~n1087;
  assign n1089 = n1088 ^ n1086;
  assign n1090 = n1089 ^ n1080;
  assign n1091 = n1090 ^ n1027;
  assign n1092 = n1082 & n1091;
  assign n1093 = n1092 ^ n1081;
  assign n1094 = n1093 ^ x103;
  assign n1095 = n1094 ^ n1071;
  assign n1096 = n1072 & n1095;
  assign n1097 = n1096 ^ n707;
  assign n1098 = n1097 ^ n608;
  assign n1099 = ~n916 & ~n1027;
  assign n1100 = n1099 ^ n920;
  assign n1101 = n1100 ^ n1097;
  assign n1102 = ~n1098 & ~n1101;
  assign n1103 = n1102 ^ n608;
  assign n1104 = n1103 ^ n514;
  assign n1105 = ~n924 & ~n1027;
  assign n1106 = n1105 ^ n942;
  assign n1107 = n1106 ^ n1103;
  assign n1108 = n1104 & ~n1107;
  assign n1109 = n1108 ^ n514;
  assign n1110 = n1109 ^ n436;
  assign n1111 = n946 & ~n1027;
  assign n1112 = n1111 ^ n949;
  assign n1113 = n1112 ^ n1109;
  assign n1114 = n1110 & ~n1113;
  assign n1115 = n1114 ^ n436;
  assign n1116 = n1115 ^ n363;
  assign n1117 = n953 & ~n1027;
  assign n1118 = n1117 ^ n956;
  assign n1119 = n1118 ^ n1115;
  assign n1120 = n1116 & ~n1119;
  assign n1121 = n1120 ^ n363;
  assign n1122 = n1121 ^ n300;
  assign n1123 = n960 & ~n1027;
  assign n1124 = n1123 ^ n963;
  assign n1125 = n1124 ^ n1121;
  assign n1126 = n1122 & n1125;
  assign n1127 = n1126 ^ n300;
  assign n1128 = n1127 ^ n243;
  assign n1129 = n967 & ~n1027;
  assign n1130 = n1129 ^ n970;
  assign n1131 = n1130 ^ n1127;
  assign n1132 = n1128 & ~n1131;
  assign n1133 = n1132 ^ n243;
  assign n1134 = n1133 ^ n210;
  assign n1135 = n974 & ~n1027;
  assign n1136 = n1135 ^ n980;
  assign n1137 = n1136 ^ n1133;
  assign n1138 = n1134 & n1137;
  assign n1139 = n1138 ^ n210;
  assign n1140 = n1139 ^ n147;
  assign n1141 = n984 & ~n1027;
  assign n1142 = n1141 ^ n987;
  assign n1143 = n1142 ^ n1139;
  assign n1144 = ~n1140 & ~n1143;
  assign n1145 = n1144 ^ n147;
  assign n1146 = n1145 ^ n132;
  assign n1147 = ~n991 & ~n1027;
  assign n1148 = n1147 ^ n997;
  assign n1149 = n1148 ^ n1145;
  assign n1150 = n1146 & ~n1149;
  assign n1151 = n1150 ^ n132;
  assign n1152 = n1151 ^ n133;
  assign n1153 = n1001 & ~n1027;
  assign n1154 = n1153 ^ n1003;
  assign n1155 = n1154 ^ n1151;
  assign n1156 = ~n1152 & ~n1155;
  assign n1157 = n1156 ^ n1151;
  assign n1158 = ~n1021 & n1157;
  assign n1159 = ~x94 & ~x95;
  assign n1160 = ~x96 & n1159;
  assign n1161 = ~n1158 & n1160;
  assign n1300 = n1158 & ~n1160;
  assign n1162 = n1146 & ~n1158;
  assign n1163 = n1162 ^ n1148;
  assign n1164 = ~n133 & n1163;
  assign n1165 = ~n1140 & ~n1158;
  assign n1166 = n1165 ^ n1142;
  assign n1167 = n1166 ^ n132;
  assign n1168 = n1027 ^ n1022;
  assign n1169 = ~n1158 & ~n1168;
  assign n1170 = n1169 ^ n1027;
  assign n1171 = n1170 ^ x100;
  assign n1172 = n1171 ^ n905;
  assign n1173 = x98 & ~x99;
  assign n1174 = ~n1158 & n1173;
  assign n1175 = ~x96 & ~x97;
  assign n1176 = ~x98 & n1175;
  assign n1177 = n1176 ^ n1027;
  assign n1178 = n1158 ^ x99;
  assign n1179 = n1178 ^ n1027;
  assign n1180 = ~n1177 & ~n1179;
  assign n1181 = n1180 ^ n1027;
  assign n1182 = ~n1174 & n1181;
  assign n1183 = n1182 ^ n1171;
  assign n1184 = ~n1172 & n1183;
  assign n1185 = n1184 ^ n905;
  assign n1186 = n1185 ^ n803;
  assign n1188 = n1027 ^ n905;
  assign n1189 = n1188 ^ n1027;
  assign n1190 = n1189 ^ n1188;
  assign n1191 = n1188 ^ n1022;
  assign n1192 = n1190 & n1191;
  assign n1193 = n1192 ^ n1188;
  assign n1194 = ~x100 & n1193;
  assign n1195 = n1194 ^ n1188;
  assign n1187 = ~x100 & ~n1027;
  assign n1196 = n1195 ^ n1187;
  assign n1197 = n1022 ^ n905;
  assign n1198 = n1197 ^ n1195;
  assign n1199 = n1195 ^ n1158;
  assign n1200 = ~n1195 & n1199;
  assign n1201 = n1200 ^ n1195;
  assign n1202 = ~n1198 & ~n1201;
  assign n1203 = n1202 ^ n1200;
  assign n1204 = n1203 ^ n1195;
  assign n1205 = n1204 ^ n1158;
  assign n1206 = n1196 & n1205;
  assign n1207 = n1206 ^ n1187;
  assign n1208 = n1207 ^ x101;
  assign n1209 = n1208 ^ n1185;
  assign n1210 = n1186 & ~n1209;
  assign n1211 = n1210 ^ n803;
  assign n1212 = n1211 ^ n707;
  assign n1221 = n908 ^ n905;
  assign n1222 = ~n1027 & ~n1221;
  assign n1223 = n1222 ^ n905;
  assign n1224 = n1223 ^ x102;
  assign n1213 = ~n1027 & n1040;
  assign n1214 = n1023 ^ n905;
  assign n1215 = n1059 ^ n1023;
  assign n1216 = ~n1214 & n1215;
  assign n1217 = n1216 ^ n1023;
  assign n1218 = ~n1213 & ~n1217;
  assign n1219 = n1218 ^ n803;
  assign n1220 = ~n1158 & n1219;
  assign n1225 = n1224 ^ n1220;
  assign n1226 = n1225 ^ n1211;
  assign n1227 = ~n1212 & n1226;
  assign n1228 = n1227 ^ n707;
  assign n1229 = n1228 ^ n608;
  assign n1230 = n1072 & ~n1158;
  assign n1231 = n1230 ^ n1094;
  assign n1232 = n1231 ^ n1228;
  assign n1233 = ~n1229 & n1232;
  assign n1234 = n1233 ^ n608;
  assign n1235 = n1234 ^ n514;
  assign n1236 = ~n1098 & ~n1158;
  assign n1237 = n1236 ^ n1100;
  assign n1238 = n1237 ^ n1234;
  assign n1239 = n1235 & n1238;
  assign n1240 = n1239 ^ n514;
  assign n1241 = n1240 ^ n436;
  assign n1242 = n1104 & ~n1158;
  assign n1243 = n1242 ^ n1106;
  assign n1244 = n1243 ^ n1240;
  assign n1245 = n1241 & ~n1244;
  assign n1246 = n1245 ^ n436;
  assign n1247 = n1246 ^ n363;
  assign n1248 = n1110 & ~n1158;
  assign n1249 = n1248 ^ n1112;
  assign n1250 = n1249 ^ n1246;
  assign n1251 = n1247 & ~n1250;
  assign n1252 = n1251 ^ n363;
  assign n1253 = n1252 ^ n300;
  assign n1254 = n1116 & ~n1158;
  assign n1255 = n1254 ^ n1118;
  assign n1256 = n1255 ^ n1252;
  assign n1257 = n1253 & ~n1256;
  assign n1258 = n1257 ^ n300;
  assign n1259 = n1258 ^ n243;
  assign n1260 = n1122 & ~n1158;
  assign n1261 = n1260 ^ n1124;
  assign n1262 = n1261 ^ n1258;
  assign n1263 = n1259 & n1262;
  assign n1264 = n1263 ^ n243;
  assign n1265 = n1264 ^ n210;
  assign n1266 = n1128 & ~n1158;
  assign n1267 = n1266 ^ n1130;
  assign n1268 = n1267 ^ n1264;
  assign n1269 = n1265 & ~n1268;
  assign n1270 = n1269 ^ n210;
  assign n1271 = n1270 ^ n147;
  assign n1272 = n1134 & ~n1158;
  assign n1273 = n1272 ^ n1136;
  assign n1274 = n1273 ^ n1270;
  assign n1275 = ~n1271 & n1274;
  assign n1276 = n1275 ^ n147;
  assign n1277 = n1276 ^ n1166;
  assign n1278 = ~n1167 & n1277;
  assign n1279 = n1278 ^ n132;
  assign n1280 = ~n1164 & ~n1279;
  assign n1281 = n1021 & ~n1151;
  assign n1282 = n132 & ~n1148;
  assign n1283 = n1145 & n1282;
  assign n1284 = ~n1021 & ~n1283;
  assign n1285 = n133 & ~n1284;
  assign n1286 = ~n1145 & ~n1148;
  assign n1287 = n129 & n133;
  assign n1288 = n1286 & n1287;
  assign n1289 = ~n1154 & ~n1288;
  assign n1290 = ~n1285 & n1289;
  assign n1291 = ~n1281 & n1290;
  assign n1292 = ~n129 & n133;
  assign n1293 = n1151 & ~n1292;
  assign n1294 = n1145 & n1148;
  assign n1295 = n133 & ~n1294;
  assign n1296 = n1154 & ~n1295;
  assign n1297 = ~n1293 & n1296;
  assign n1298 = ~n1291 & ~n1297;
  assign n1299 = ~n1280 & ~n1298;
  assign n1301 = n1300 ^ n1299;
  assign n1302 = n1301 ^ x97;
  assign n1303 = n1302 ^ n1299;
  assign n1304 = n1303 ^ n1301;
  assign n1305 = ~x96 & ~n1299;
  assign n1306 = n1305 ^ n1301;
  assign n1307 = ~n1304 & ~n1306;
  assign n1308 = n1307 ^ n1302;
  assign n1309 = ~n1161 & ~n1308;
  assign n1310 = n1309 ^ n1027;
  assign n1311 = n1175 ^ n1158;
  assign n1312 = ~n1299 & ~n1311;
  assign n1313 = n1312 ^ n1158;
  assign n1314 = n1313 ^ x98;
  assign n1315 = n1314 ^ n1309;
  assign n1316 = n1310 & n1315;
  assign n1317 = n1316 ^ n1027;
  assign n1318 = n1317 ^ n905;
  assign n1320 = n1158 ^ n1027;
  assign n1321 = n1320 ^ n1158;
  assign n1322 = n1321 ^ n1320;
  assign n1323 = n1320 ^ n1175;
  assign n1324 = n1322 & n1323;
  assign n1325 = n1324 ^ n1320;
  assign n1326 = ~x98 & n1325;
  assign n1327 = n1326 ^ n1320;
  assign n1319 = ~x98 & ~n1158;
  assign n1328 = n1327 ^ n1319;
  assign n1329 = n1175 ^ n1027;
  assign n1330 = n1329 ^ n1327;
  assign n1331 = n1327 ^ n1299;
  assign n1332 = ~n1327 & n1331;
  assign n1333 = n1332 ^ n1327;
  assign n1334 = ~n1330 & ~n1333;
  assign n1335 = n1334 ^ n1332;
  assign n1336 = n1335 ^ n1327;
  assign n1337 = n1336 ^ n1299;
  assign n1338 = n1328 & n1337;
  assign n1339 = n1338 ^ n1319;
  assign n1340 = n1339 ^ x99;
  assign n1341 = n1340 ^ n1317;
  assign n1342 = n1318 & ~n1341;
  assign n1343 = n1342 ^ n905;
  assign n1344 = n1343 ^ n803;
  assign n1345 = n1182 ^ n905;
  assign n1346 = ~n1299 & n1345;
  assign n1347 = n1346 ^ n1171;
  assign n1348 = n1347 ^ n1343;
  assign n1349 = n1344 & n1348;
  assign n1350 = n1349 ^ n803;
  assign n1351 = n1350 ^ n707;
  assign n1352 = n1186 & ~n1299;
  assign n1353 = n1352 ^ n1208;
  assign n1354 = n1353 ^ n1350;
  assign n1355 = ~n1351 & ~n1354;
  assign n1356 = n1355 ^ n707;
  assign n1357 = n1356 ^ n608;
  assign n1358 = ~n1212 & ~n1299;
  assign n1359 = n1358 ^ n1225;
  assign n1360 = n1359 ^ n1356;
  assign n1361 = ~n1357 & ~n1360;
  assign n1362 = n1361 ^ n608;
  assign n1363 = n1362 ^ n514;
  assign n1364 = ~n1229 & ~n1299;
  assign n1365 = n1364 ^ n1231;
  assign n1366 = n1365 ^ n1362;
  assign n1367 = n1363 & ~n1366;
  assign n1368 = n1367 ^ n514;
  assign n1369 = n1368 ^ n436;
  assign n1370 = ~n1271 & ~n1299;
  assign n1371 = n1370 ^ n1273;
  assign n1372 = n1265 & ~n1299;
  assign n1373 = n1372 ^ n1267;
  assign n1374 = n1373 ^ n147;
  assign n1375 = n1259 & ~n1299;
  assign n1376 = n1375 ^ n1261;
  assign n1377 = n1376 ^ n210;
  assign n1378 = n1235 & ~n1299;
  assign n1379 = n1378 ^ n1237;
  assign n1380 = n1379 ^ n1368;
  assign n1381 = n1369 & n1380;
  assign n1382 = n1381 ^ n436;
  assign n1383 = n1382 ^ n363;
  assign n1384 = n1241 & ~n1299;
  assign n1385 = n1384 ^ n1243;
  assign n1386 = n1385 ^ n1382;
  assign n1387 = n1383 & ~n1386;
  assign n1388 = n1387 ^ n363;
  assign n1389 = n1388 ^ n300;
  assign n1390 = n1247 & ~n1299;
  assign n1391 = n1390 ^ n1249;
  assign n1392 = n1391 ^ n1388;
  assign n1393 = n1389 & ~n1392;
  assign n1394 = n1393 ^ n300;
  assign n1395 = n1394 ^ n243;
  assign n1396 = n1253 & ~n1299;
  assign n1397 = n1396 ^ n1255;
  assign n1398 = n1397 ^ n1394;
  assign n1399 = n1395 & ~n1398;
  assign n1400 = n1399 ^ n243;
  assign n1401 = n1400 ^ n1376;
  assign n1402 = ~n1377 & n1401;
  assign n1403 = n1402 ^ n210;
  assign n1404 = n1403 ^ n1373;
  assign n1405 = ~n1374 & ~n1404;
  assign n1406 = n1405 ^ n147;
  assign n1407 = ~n1371 & ~n1406;
  assign n1408 = ~n1166 & n1299;
  assign n1409 = n1276 ^ n1167;
  assign n1410 = n1299 ^ n1276;
  assign n1411 = n1277 ^ n1276;
  assign n1412 = n1410 & n1411;
  assign n1413 = n1412 ^ n1276;
  assign n1414 = ~n1409 & ~n1413;
  assign n1415 = ~n1408 & ~n1414;
  assign n1416 = n1279 ^ n1163;
  assign n1417 = n1416 ^ n1163;
  assign n1418 = n1163 & n1298;
  assign n1419 = n1418 ^ n1163;
  assign n1420 = ~n1417 & ~n1419;
  assign n1421 = n1420 ^ n1163;
  assign n1422 = ~n133 & n1421;
  assign n1423 = ~n1415 & n1422;
  assign n1424 = ~n1166 & n1276;
  assign n1425 = n1422 & n1424;
  assign n1426 = ~n1423 & ~n1425;
  assign n1427 = n1407 & n1426;
  assign n1428 = ~n132 & ~n1423;
  assign n1429 = ~n1406 & n1428;
  assign n1430 = n1163 & n1414;
  assign n1431 = n1166 & ~n1276;
  assign n1432 = n132 & n1431;
  assign n1433 = ~n1299 & n1432;
  assign n1434 = ~n1371 & ~n1433;
  assign n1435 = n1430 & ~n1434;
  assign n1437 = ~n1166 & ~n1298;
  assign n1436 = n132 & ~n1418;
  assign n1438 = n1437 ^ n1436;
  assign n1439 = n1437 ^ n1424;
  assign n1440 = n1439 ^ n1424;
  assign n1441 = ~n147 & n1270;
  assign n1442 = n1273 & ~n1441;
  assign n1443 = n1442 ^ n1424;
  assign n1444 = n1440 & ~n1443;
  assign n1445 = n1444 ^ n1424;
  assign n1446 = n1438 & ~n1445;
  assign n1447 = n1446 ^ n1436;
  assign n1448 = ~n1435 & ~n1447;
  assign n1449 = n1448 ^ n1421;
  assign n1450 = n133 & ~n1449;
  assign n1451 = n1450 ^ n1421;
  assign n1452 = ~n1429 & n1451;
  assign n1453 = ~n1427 & n1452;
  assign n1454 = ~n132 & ~n1371;
  assign n1455 = n1276 & ~n1299;
  assign n1456 = n1455 ^ n1166;
  assign n1457 = n1454 & n1456;
  assign n1458 = n1453 & ~n1457;
  assign n1459 = n1369 & ~n1458;
  assign n1460 = n1459 ^ n1379;
  assign n1461 = n1460 ^ n363;
  assign n1462 = n1363 & ~n1458;
  assign n1463 = n1462 ^ n1365;
  assign n1464 = n1463 ^ n436;
  assign n1465 = ~n1357 & ~n1458;
  assign n1466 = n1465 ^ n1359;
  assign n1467 = n514 & ~n1466;
  assign n1468 = n1467 ^ n1463;
  assign n1469 = n1464 & n1468;
  assign n1470 = n1469 ^ n1463;
  assign n1471 = n1470 ^ n1460;
  assign n1472 = n1471 ^ n1460;
  assign n1473 = ~n436 & ~n1463;
  assign n1474 = ~n514 & n1466;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~x92 & ~x93;
  assign n1477 = ~n1299 & n1476;
  assign n1478 = ~x94 & n1477;
  assign n1479 = n1458 ^ x95;
  assign n1480 = x94 & n1299;
  assign n1481 = n1299 & ~n1476;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = n1482 ^ x94;
  assign n1484 = n1483 ^ n1482;
  assign n1485 = n1482 ^ n1458;
  assign n1486 = n1485 ^ n1482;
  assign n1487 = n1484 & ~n1486;
  assign n1488 = n1487 ^ n1482;
  assign n1489 = ~n1479 & n1488;
  assign n1490 = n1489 ^ n1482;
  assign n1491 = ~n1478 & ~n1490;
  assign n1492 = n1491 ^ n1158;
  assign n1493 = n1299 ^ n1159;
  assign n1494 = ~n1458 & ~n1493;
  assign n1495 = n1494 ^ n1299;
  assign n1496 = n1495 ^ x96;
  assign n1497 = n1496 ^ n1491;
  assign n1498 = n1492 & n1497;
  assign n1499 = n1498 ^ n1158;
  assign n1500 = n1499 ^ n1027;
  assign n1502 = x96 & n1158;
  assign n1501 = n1160 ^ n1158;
  assign n1503 = n1502 ^ n1501;
  assign n1504 = ~n1299 & ~n1503;
  assign n1505 = n1504 ^ n1501;
  assign n1506 = n1505 ^ n1305;
  assign n1507 = n1159 ^ n1158;
  assign n1508 = n1507 ^ n1505;
  assign n1509 = n1505 ^ n1458;
  assign n1510 = n1505 & ~n1509;
  assign n1511 = n1510 ^ n1505;
  assign n1512 = n1508 & n1511;
  assign n1513 = n1512 ^ n1510;
  assign n1514 = n1513 ^ n1505;
  assign n1515 = n1514 ^ n1458;
  assign n1516 = ~n1506 & ~n1515;
  assign n1517 = n1516 ^ n1305;
  assign n1518 = n1517 ^ x97;
  assign n1519 = n1518 ^ n1499;
  assign n1520 = n1500 & ~n1519;
  assign n1521 = n1520 ^ n1027;
  assign n1522 = n1521 ^ n905;
  assign n1523 = n1310 & ~n1458;
  assign n1524 = n1523 ^ n1314;
  assign n1525 = n1524 ^ n1521;
  assign n1526 = n1522 & n1525;
  assign n1527 = n1526 ^ n905;
  assign n1528 = n1527 ^ n803;
  assign n1529 = n1318 & ~n1458;
  assign n1530 = n1529 ^ n1340;
  assign n1531 = n1530 ^ n1527;
  assign n1532 = n1528 & ~n1531;
  assign n1533 = n1532 ^ n803;
  assign n1534 = n1533 ^ n707;
  assign n1535 = n1344 & ~n1458;
  assign n1536 = n1535 ^ n1347;
  assign n1537 = n1536 ^ n1533;
  assign n1538 = ~n1534 & n1537;
  assign n1539 = n1538 ^ n707;
  assign n1540 = n1539 ^ n608;
  assign n1541 = ~n1351 & ~n1458;
  assign n1542 = n1541 ^ n1353;
  assign n1543 = n1542 ^ n1539;
  assign n1544 = ~n1540 & n1543;
  assign n1545 = n1544 ^ n608;
  assign n1546 = n1475 & n1545;
  assign n1547 = n1546 ^ n1460;
  assign n1548 = n1547 ^ n1460;
  assign n1549 = ~n1472 & ~n1548;
  assign n1550 = n1549 ^ n1460;
  assign n1551 = ~n1461 & ~n1550;
  assign n1552 = n1551 ^ n363;
  assign n1553 = n1552 ^ n300;
  assign n1554 = n1383 & ~n1458;
  assign n1555 = n1554 ^ n1385;
  assign n1556 = n1555 ^ n1552;
  assign n1557 = n1553 & ~n1556;
  assign n1558 = n1557 ^ n300;
  assign n1559 = n1558 ^ n243;
  assign n1560 = n1389 & ~n1458;
  assign n1561 = n1560 ^ n1391;
  assign n1562 = n1561 ^ n1558;
  assign n1563 = n1559 & ~n1562;
  assign n1564 = n1563 ^ n243;
  assign n1565 = n1564 ^ n210;
  assign n1566 = n1395 & ~n1458;
  assign n1567 = n1566 ^ n1397;
  assign n1568 = n1567 ^ n1564;
  assign n1569 = n1565 & ~n1568;
  assign n1570 = n1569 ^ n210;
  assign n1571 = n1570 ^ n147;
  assign n1572 = n1406 ^ n132;
  assign n1573 = ~n1458 & n1572;
  assign n1574 = n1573 ^ n1371;
  assign n1575 = ~n133 & n1574;
  assign n1576 = n1400 ^ n210;
  assign n1577 = ~n1458 & n1576;
  assign n1578 = n1577 ^ n1376;
  assign n1579 = n1578 ^ n1570;
  assign n1580 = ~n1571 & n1579;
  assign n1581 = n1580 ^ n147;
  assign n1582 = n1581 ^ n132;
  assign n1583 = n1403 ^ n147;
  assign n1584 = ~n1458 & ~n1583;
  assign n1585 = n1584 ^ n1373;
  assign n1586 = n1585 ^ n1581;
  assign n1587 = n1582 & n1586;
  assign n1588 = n1587 ^ n132;
  assign n1589 = ~n1575 & ~n1588;
  assign n1590 = n1276 ^ n132;
  assign n1591 = ~n1299 & n1590;
  assign n1592 = n1591 ^ n1166;
  assign n1595 = n1371 & n1406;
  assign n1596 = n1292 & ~n1451;
  assign n1597 = n1595 & n1596;
  assign n1598 = n1592 & ~n1597;
  assign n1593 = n1371 & n1452;
  assign n1594 = ~n1592 & ~n1593;
  assign n1599 = n1598 ^ n1594;
  assign n1600 = ~n1371 & n1458;
  assign n1601 = ~n132 & ~n1595;
  assign n1602 = ~n1407 & n1601;
  assign n1603 = ~n1600 & n1602;
  assign n1604 = n132 & n1407;
  assign n1605 = ~n1453 & n1604;
  assign n1606 = n133 & ~n1605;
  assign n1607 = ~n1603 & n1606;
  assign n1608 = n1607 ^ n1598;
  assign n1609 = ~n1407 & ~n1601;
  assign n1610 = ~n133 & ~n1609;
  assign n1611 = ~n1458 & n1610;
  assign n1612 = n1611 ^ n1598;
  assign n1613 = ~n1598 & n1612;
  assign n1614 = n1613 ^ n1598;
  assign n1615 = ~n1608 & ~n1614;
  assign n1616 = n1615 ^ n1613;
  assign n1617 = n1616 ^ n1598;
  assign n1618 = n1617 ^ n1611;
  assign n1619 = n1599 & n1618;
  assign n1620 = n1619 ^ n1594;
  assign n1621 = ~n1589 & ~n1620;
  assign n1622 = ~n1571 & ~n1621;
  assign n1623 = n1622 ^ n1578;
  assign n1624 = n1545 ^ n514;
  assign n1625 = ~n1621 & n1624;
  assign n1626 = n1625 ^ n1466;
  assign n1627 = n1626 ^ n436;
  assign n1628 = ~n1540 & ~n1621;
  assign n1629 = n1628 ^ n1542;
  assign n1630 = n1629 ^ n514;
  assign n1631 = ~n1534 & ~n1621;
  assign n1632 = n1631 ^ n1536;
  assign n1633 = ~n608 & n1632;
  assign n1634 = n1633 ^ n1629;
  assign n1635 = n1630 & ~n1634;
  assign n1636 = n1635 ^ n1629;
  assign n1637 = n1636 ^ n1626;
  assign n1638 = n1637 ^ n1626;
  assign n1639 = n608 & ~n1632;
  assign n1640 = n514 & n1629;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = n1522 & ~n1621;
  assign n1643 = n1642 ^ n1524;
  assign n1644 = n1643 ^ n803;
  assign n1645 = n1500 & ~n1621;
  assign n1646 = n1645 ^ n1518;
  assign n1647 = n1646 ^ n905;
  assign n1648 = n1492 & ~n1621;
  assign n1649 = n1648 ^ n1496;
  assign n1650 = n1027 & ~n1649;
  assign n1651 = n1650 ^ n1646;
  assign n1652 = n1647 & n1651;
  assign n1653 = n1652 ^ n1646;
  assign n1654 = n1653 ^ n1643;
  assign n1655 = n1654 ^ n1643;
  assign n1656 = ~n905 & ~n1646;
  assign n1657 = ~n1027 & n1649;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = n1476 ^ n1458;
  assign n1660 = ~n1621 & ~n1659;
  assign n1661 = n1660 ^ n1458;
  assign n1662 = n1661 ^ x94;
  assign n1663 = n1662 ^ n1299;
  assign n1664 = ~x90 & ~x91;
  assign n1665 = ~n1458 & n1664;
  assign n1666 = ~x92 & n1665;
  assign n1667 = x92 & n1458;
  assign n1668 = n1458 & ~n1664;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n1669 ^ n1621;
  assign n1671 = n1670 ^ x93;
  assign n1672 = n1671 ^ n1621;
  assign n1673 = n1672 ^ n1670;
  assign n1674 = ~x92 & ~n1621;
  assign n1675 = n1674 ^ n1670;
  assign n1676 = ~n1673 & n1675;
  assign n1677 = n1676 ^ n1671;
  assign n1678 = ~n1666 & n1677;
  assign n1679 = n1678 ^ n1662;
  assign n1680 = ~n1663 & n1679;
  assign n1681 = n1680 ^ n1299;
  assign n1682 = n1681 ^ n1158;
  assign n1684 = n1480 ^ n1478;
  assign n1685 = n1684 ^ n1480;
  assign n1686 = n1482 ^ n1480;
  assign n1687 = n1686 ^ n1480;
  assign n1688 = ~n1685 & n1687;
  assign n1689 = n1688 ^ n1480;
  assign n1690 = n1458 & n1689;
  assign n1691 = n1690 ^ n1480;
  assign n1683 = ~x94 & ~n1458;
  assign n1692 = n1691 ^ n1683;
  assign n1693 = n1476 ^ n1299;
  assign n1694 = n1693 ^ n1691;
  assign n1695 = n1691 ^ n1621;
  assign n1696 = ~n1691 & n1695;
  assign n1697 = n1696 ^ n1691;
  assign n1698 = ~n1694 & ~n1697;
  assign n1699 = n1698 ^ n1696;
  assign n1700 = n1699 ^ n1691;
  assign n1701 = n1700 ^ n1621;
  assign n1702 = n1692 & n1701;
  assign n1703 = n1702 ^ n1683;
  assign n1704 = n1703 ^ x95;
  assign n1705 = n1704 ^ n1681;
  assign n1706 = n1682 & ~n1705;
  assign n1707 = n1706 ^ n1158;
  assign n1708 = n1658 & n1707;
  assign n1709 = n1708 ^ n1643;
  assign n1710 = n1709 ^ n1643;
  assign n1711 = ~n1655 & ~n1710;
  assign n1712 = n1711 ^ n1643;
  assign n1713 = ~n1644 & ~n1712;
  assign n1714 = n1713 ^ n803;
  assign n1715 = n1714 ^ n707;
  assign n1716 = n1528 & ~n1621;
  assign n1717 = n1716 ^ n1530;
  assign n1718 = n1717 ^ n1714;
  assign n1719 = ~n1715 & ~n1718;
  assign n1720 = n1719 ^ n707;
  assign n1721 = n1641 & n1720;
  assign n1722 = n1721 ^ n1626;
  assign n1723 = n1722 ^ n1626;
  assign n1724 = n1638 & ~n1723;
  assign n1725 = n1724 ^ n1626;
  assign n1726 = ~n1627 & n1725;
  assign n1727 = n1726 ^ n436;
  assign n1728 = n1727 ^ n363;
  assign n1729 = n1466 ^ n514;
  assign n1730 = n1545 ^ n1466;
  assign n1731 = ~n1729 & n1730;
  assign n1732 = n1731 ^ n514;
  assign n1733 = n1732 ^ n436;
  assign n1734 = ~n1621 & n1733;
  assign n1735 = n1734 ^ n1463;
  assign n1736 = n1735 ^ n1727;
  assign n1737 = n1728 & ~n1736;
  assign n1738 = n1737 ^ n363;
  assign n1739 = n1738 ^ n300;
  assign n1740 = n1732 ^ n1463;
  assign n1741 = n1464 & ~n1740;
  assign n1742 = n1741 ^ n436;
  assign n1743 = n1742 ^ n363;
  assign n1744 = ~n1621 & n1743;
  assign n1745 = n1744 ^ n1460;
  assign n1746 = n1745 ^ n1738;
  assign n1747 = n1739 & n1746;
  assign n1748 = n1747 ^ n300;
  assign n1749 = n1748 ^ n243;
  assign n1750 = n1553 & ~n1621;
  assign n1751 = n1750 ^ n1555;
  assign n1752 = n1751 ^ n1748;
  assign n1753 = n1749 & ~n1752;
  assign n1754 = n1753 ^ n243;
  assign n1755 = n1754 ^ n210;
  assign n1756 = n1559 & ~n1621;
  assign n1757 = n1756 ^ n1561;
  assign n1758 = n1757 ^ n1754;
  assign n1759 = n1755 & ~n1758;
  assign n1760 = n1759 ^ n210;
  assign n1761 = n1760 ^ n147;
  assign n1762 = n1565 & ~n1621;
  assign n1763 = n1762 ^ n1567;
  assign n1764 = n1763 ^ n1760;
  assign n1765 = ~n1761 & ~n1764;
  assign n1766 = n1765 ^ n147;
  assign n1767 = ~n1623 & ~n1766;
  assign n1768 = n132 & ~n1767;
  assign n1769 = n1623 & n1766;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = n133 & ~n1766;
  assign n1772 = n132 & n1581;
  assign n1773 = ~n132 & ~n1581;
  assign n1774 = ~n1621 & ~n1773;
  assign n1775 = ~n1772 & n1774;
  assign n1776 = n1775 ^ n1585;
  assign n1777 = ~n1771 & ~n1776;
  assign n1778 = n1770 & ~n1777;
  assign n1779 = ~n132 & n1623;
  assign n1780 = ~n1581 & n1585;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = n1774 ^ n1581;
  assign n1783 = n1585 & ~n1782;
  assign n1784 = n1783 ^ n1581;
  assign n1785 = n1574 & ~n1784;
  assign n1786 = ~n1781 & n1785;
  assign n1787 = ~n147 & n1570;
  assign n1788 = n1578 & ~n1787;
  assign n1789 = ~n132 & ~n1788;
  assign n1790 = n1621 & ~n1789;
  assign n1791 = ~n1574 & n1772;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n1585 & ~n1792;
  assign n1794 = n133 & ~n1793;
  assign n1795 = ~n1786 & n1794;
  assign n1796 = n1588 ^ n1574;
  assign n1797 = n1574 ^ n133;
  assign n1798 = n1620 ^ n133;
  assign n1799 = n1798 ^ n133;
  assign n1800 = n1797 & ~n1799;
  assign n1801 = n1800 ^ n133;
  assign n1802 = n1796 & ~n1801;
  assign n1803 = ~n1795 & ~n1802;
  assign n1804 = ~n1778 & n1803;
  assign n1805 = n1766 ^ n132;
  assign n1806 = ~n1804 & n1805;
  assign n1807 = n1806 ^ n1623;
  assign n1808 = ~n1761 & ~n1804;
  assign n1809 = n1808 ^ n1763;
  assign n1815 = n132 & n1809;
  assign n1816 = ~n1715 & ~n1804;
  assign n1817 = n1816 ^ n1717;
  assign n1818 = ~n608 & ~n1817;
  assign n1819 = n1720 ^ n608;
  assign n1820 = ~n1804 & ~n1819;
  assign n1821 = n1820 ^ n1632;
  assign n1822 = ~n514 & n1821;
  assign n1823 = ~n1818 & ~n1822;
  assign n1824 = n1649 ^ n1027;
  assign n1825 = n1707 ^ n1649;
  assign n1826 = ~n1824 & n1825;
  assign n1827 = n1826 ^ n1027;
  assign n1828 = n1827 ^ n905;
  assign n1829 = ~n1804 & n1828;
  assign n1830 = n1829 ^ n1646;
  assign n1831 = n1830 ^ n803;
  assign n1832 = n1707 ^ n1027;
  assign n1833 = ~n1804 & n1832;
  assign n1834 = n1833 ^ n1649;
  assign n1835 = n1834 ^ n905;
  assign n1836 = ~x88 & ~x89;
  assign n1837 = ~n1621 & n1836;
  assign n1838 = ~x90 & n1837;
  assign n1839 = n1804 ^ x91;
  assign n1840 = x90 & n1621;
  assign n1841 = n1621 & ~n1836;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = n1842 ^ x90;
  assign n1844 = n1843 ^ n1842;
  assign n1845 = n1842 ^ n1804;
  assign n1846 = n1845 ^ n1842;
  assign n1847 = n1844 & ~n1846;
  assign n1848 = n1847 ^ n1842;
  assign n1849 = ~n1839 & n1848;
  assign n1850 = n1849 ^ n1842;
  assign n1851 = ~n1838 & ~n1850;
  assign n1852 = n1851 ^ n1458;
  assign n1853 = n1664 ^ n1621;
  assign n1854 = ~n1804 & ~n1853;
  assign n1855 = n1854 ^ n1621;
  assign n1856 = n1855 ^ x92;
  assign n1857 = n1856 ^ n1851;
  assign n1858 = n1852 & n1857;
  assign n1859 = n1858 ^ n1458;
  assign n1860 = n1859 ^ n1299;
  assign n1861 = ~n1666 & n1669;
  assign n1862 = n1861 ^ n1667;
  assign n1863 = n1621 & n1862;
  assign n1864 = n1863 ^ n1667;
  assign n1865 = n1864 ^ n1674;
  assign n1866 = n1664 ^ n1458;
  assign n1867 = n1866 ^ n1864;
  assign n1868 = n1864 ^ n1804;
  assign n1869 = ~n1864 & n1868;
  assign n1870 = n1869 ^ n1864;
  assign n1871 = ~n1867 & ~n1870;
  assign n1872 = n1871 ^ n1869;
  assign n1873 = n1872 ^ n1864;
  assign n1874 = n1873 ^ n1804;
  assign n1875 = n1865 & n1874;
  assign n1876 = n1875 ^ n1674;
  assign n1877 = n1876 ^ x93;
  assign n1878 = n1877 ^ n1859;
  assign n1879 = n1860 & ~n1878;
  assign n1880 = n1879 ^ n1299;
  assign n1881 = n1880 ^ n1158;
  assign n1882 = n1678 ^ n1299;
  assign n1883 = ~n1804 & n1882;
  assign n1884 = n1883 ^ n1662;
  assign n1885 = n1884 ^ n1880;
  assign n1886 = n1881 & n1885;
  assign n1887 = n1886 ^ n1158;
  assign n1888 = n1887 ^ n1027;
  assign n1889 = n1682 & ~n1804;
  assign n1890 = n1889 ^ n1704;
  assign n1891 = n1890 ^ n1887;
  assign n1892 = n1888 & ~n1891;
  assign n1893 = n1892 ^ n1027;
  assign n1894 = n1893 ^ n1834;
  assign n1895 = ~n1835 & n1894;
  assign n1896 = n1895 ^ n905;
  assign n1897 = n1896 ^ n1830;
  assign n1898 = n1831 & ~n1897;
  assign n1899 = n1898 ^ n803;
  assign n1900 = n1899 ^ n707;
  assign n1901 = n1827 ^ n1646;
  assign n1902 = n1647 & ~n1901;
  assign n1903 = n1902 ^ n905;
  assign n1904 = n1903 ^ n803;
  assign n1905 = ~n1804 & n1904;
  assign n1906 = n1905 ^ n1643;
  assign n1907 = n1906 ^ n1899;
  assign n1908 = ~n1900 & n1907;
  assign n1909 = n1908 ^ n707;
  assign n1910 = n1823 & ~n1909;
  assign n1911 = n1821 ^ n514;
  assign n1912 = n608 & n1817;
  assign n1913 = n1912 ^ n1821;
  assign n1914 = ~n1911 & n1913;
  assign n1915 = n1914 ^ n514;
  assign n1916 = ~n1910 & ~n1915;
  assign n1917 = n1916 ^ n436;
  assign n1918 = n1632 ^ n608;
  assign n1919 = n1720 ^ n1632;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = n1920 ^ n608;
  assign n1922 = n1921 ^ n514;
  assign n1923 = ~n1804 & n1922;
  assign n1924 = n1923 ^ n1629;
  assign n1925 = n1924 ^ n1916;
  assign n1926 = ~n1917 & n1925;
  assign n1927 = n1926 ^ n436;
  assign n1928 = n1927 ^ n363;
  assign n1929 = n1921 ^ n1629;
  assign n1930 = n1630 & ~n1929;
  assign n1931 = n1930 ^ n514;
  assign n1932 = n1931 ^ n436;
  assign n1933 = ~n1804 & n1932;
  assign n1934 = n1933 ^ n1626;
  assign n1935 = n1934 ^ n1927;
  assign n1936 = n1928 & n1935;
  assign n1937 = n1936 ^ n363;
  assign n1938 = n1937 ^ n300;
  assign n1939 = n1728 & ~n1804;
  assign n1940 = n1939 ^ n1735;
  assign n1941 = n1940 ^ n1937;
  assign n1942 = n1938 & ~n1941;
  assign n1943 = n1942 ^ n300;
  assign n1944 = n1943 ^ n243;
  assign n1945 = n1739 & ~n1804;
  assign n1946 = n1945 ^ n1745;
  assign n1947 = n1946 ^ n1943;
  assign n1948 = n1944 & n1947;
  assign n1949 = n1948 ^ n243;
  assign n1950 = n1949 ^ n210;
  assign n1951 = n1749 & ~n1804;
  assign n1952 = n1951 ^ n1751;
  assign n1953 = n1952 ^ n1949;
  assign n1954 = n1950 & ~n1953;
  assign n1955 = n1954 ^ n210;
  assign n1956 = n1955 ^ n147;
  assign n1810 = n1755 & ~n1804;
  assign n1811 = n1810 ^ n1757;
  assign n1957 = n1955 ^ n1811;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = n1958 ^ n147;
  assign n1960 = n1815 & ~n1959;
  assign n1961 = ~n147 & n1955;
  assign n1812 = ~n1809 & ~n1811;
  assign n1962 = ~n132 & ~n1812;
  assign n1963 = ~n1961 & n1962;
  assign n1964 = n1811 ^ n1809;
  assign n1965 = n147 & ~n1955;
  assign n1966 = n1965 ^ n1809;
  assign n1967 = n1966 ^ n1809;
  assign n1968 = n1964 & n1967;
  assign n1969 = n1968 ^ n1809;
  assign n1970 = n1963 & ~n1969;
  assign n1971 = ~n1960 & ~n1970;
  assign n1813 = n132 & ~n1809;
  assign n1814 = ~n1812 & ~n1813;
  assign n1972 = n1971 ^ n1814;
  assign n1973 = ~n132 & ~n147;
  assign n1974 = n1955 & n1973;
  assign n1975 = n1974 ^ n1971;
  assign n1976 = ~n132 & n1809;
  assign n1977 = n1959 & ~n1976;
  assign n1978 = ~n133 & n1807;
  assign n1979 = ~n1813 & ~n1978;
  assign n1980 = ~n1977 & n1979;
  assign n1981 = n1766 ^ n1623;
  assign n1982 = n1981 ^ n1766;
  assign n1983 = n1803 ^ n1766;
  assign n1984 = ~n1982 & n1983;
  assign n1985 = n1984 ^ n1766;
  assign n1986 = ~n1776 & ~n1985;
  assign n1987 = ~n1767 & n1986;
  assign n1988 = n1287 & ~n1987;
  assign n1989 = ~n1768 & ~n1776;
  assign n1990 = n1776 & ~n1803;
  assign n1991 = n1769 & n1990;
  assign n1992 = n133 & ~n1991;
  assign n1993 = ~n1989 & n1992;
  assign n1994 = ~n1988 & ~n1993;
  assign n1995 = n132 & n1766;
  assign n1996 = ~n1776 & ~n1803;
  assign n1997 = ~n1623 & ~n1996;
  assign n1998 = ~n1995 & n1997;
  assign n1999 = ~n133 & ~n1998;
  assign n2000 = n1776 ^ n1770;
  assign n2001 = n2000 ^ n1770;
  assign n2002 = ~n132 & ~n1766;
  assign n2003 = n2002 ^ n1770;
  assign n2004 = n2001 & ~n2003;
  assign n2005 = n2004 ^ n1770;
  assign n2006 = n1999 & n2005;
  assign n2007 = n1994 & ~n2006;
  assign n2008 = n1623 & ~n1776;
  assign n2009 = n1803 & n2008;
  assign n2010 = ~n2007 & ~n2009;
  assign n2011 = ~n1980 & ~n2010;
  assign n2012 = n2011 ^ n1971;
  assign n2013 = n1971 & ~n2012;
  assign n2014 = n2013 ^ n1971;
  assign n2015 = n1975 & n2014;
  assign n2016 = n2015 ^ n2013;
  assign n2017 = n2016 ^ n1971;
  assign n2018 = n2017 ^ n2011;
  assign n2019 = n1972 & ~n2018;
  assign n2020 = n2019 ^ n1814;
  assign n2021 = n1807 & ~n2020;
  assign n2022 = ~n1807 & n2010;
  assign n2023 = n1813 & n2022;
  assign n2024 = n1959 & n2023;
  assign n2025 = ~n2021 & ~n2024;
  assign n2026 = n133 & ~n2025;
  assign n2027 = ~n1813 & ~n1977;
  assign n2028 = n2027 ^ n1807;
  assign n2029 = n2027 ^ n2010;
  assign n2030 = n2027 ^ n133;
  assign n2031 = n2027 & ~n2030;
  assign n2032 = n2031 ^ n2027;
  assign n2033 = ~n2029 & n2032;
  assign n2034 = n2033 ^ n2031;
  assign n2035 = n2034 ^ n2027;
  assign n2036 = n2035 ^ n133;
  assign n2037 = ~n2028 & ~n2036;
  assign n2038 = n2037 ^ n133;
  assign n2039 = ~n2026 & n2038;
  assign n2040 = ~n1956 & ~n2011;
  assign n2041 = n2040 ^ n1811;
  assign n2042 = ~n132 & n2041;
  assign n2043 = n1959 ^ n132;
  assign n2044 = ~n2011 & n2043;
  assign n2045 = n2044 ^ n1809;
  assign n2046 = n2042 & n2045;
  assign n2047 = ~n2039 & ~n2046;
  assign n2048 = n1928 & ~n2011;
  assign n2049 = n2048 ^ n1934;
  assign n2050 = n2049 ^ n300;
  assign n2051 = ~n1917 & ~n2011;
  assign n2052 = n2051 ^ n1924;
  assign n2053 = n2052 ^ n363;
  assign n2054 = n1860 & ~n2011;
  assign n2055 = n2054 ^ n1877;
  assign n2056 = n2055 ^ n1158;
  assign n2057 = n1852 & ~n2011;
  assign n2058 = n2057 ^ n1856;
  assign n2059 = n2058 ^ n1299;
  assign n2061 = n1840 ^ n1838;
  assign n2062 = n2061 ^ n1840;
  assign n2063 = n1842 ^ n1840;
  assign n2064 = n2063 ^ n1840;
  assign n2065 = ~n2062 & n2064;
  assign n2066 = n2065 ^ n1840;
  assign n2067 = n1804 & n2066;
  assign n2068 = n2067 ^ n1840;
  assign n2060 = ~x90 & ~n1804;
  assign n2069 = n2068 ^ n2060;
  assign n2070 = n1836 ^ n1621;
  assign n2071 = n2070 ^ n2068;
  assign n2072 = n2068 ^ n2011;
  assign n2073 = ~n2068 & n2072;
  assign n2074 = n2073 ^ n2068;
  assign n2075 = ~n2071 & ~n2074;
  assign n2076 = n2075 ^ n2073;
  assign n2077 = n2076 ^ n2068;
  assign n2078 = n2077 ^ n2011;
  assign n2079 = n2069 & n2078;
  assign n2080 = n2079 ^ n2060;
  assign n2081 = n2080 ^ x91;
  assign n2082 = n2081 ^ n1458;
  assign n2083 = ~x86 & ~x87;
  assign n2084 = ~n1804 & n2083;
  assign n2085 = ~x88 & n2084;
  assign n2086 = n2011 ^ x89;
  assign n2087 = x88 & n1804;
  assign n2088 = n1804 & ~n2083;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = n2089 ^ x88;
  assign n2091 = n2090 ^ n2089;
  assign n2092 = n2089 ^ n2011;
  assign n2093 = n2092 ^ n2089;
  assign n2094 = n2091 & ~n2093;
  assign n2095 = n2094 ^ n2089;
  assign n2096 = ~n2086 & n2095;
  assign n2097 = n2096 ^ n2089;
  assign n2098 = ~n2085 & ~n2097;
  assign n2099 = n2098 ^ n1621;
  assign n2100 = n1836 ^ n1804;
  assign n2101 = ~n2011 & ~n2100;
  assign n2102 = n2101 ^ n1804;
  assign n2103 = n2102 ^ x90;
  assign n2104 = n2103 ^ n2098;
  assign n2105 = n2099 & n2104;
  assign n2106 = n2105 ^ n1621;
  assign n2107 = n2106 ^ n2081;
  assign n2108 = n2082 & ~n2107;
  assign n2109 = n2108 ^ n1458;
  assign n2110 = n2109 ^ n2058;
  assign n2111 = ~n2059 & n2110;
  assign n2112 = n2111 ^ n1299;
  assign n2113 = n2112 ^ n2055;
  assign n2114 = n2056 & ~n2113;
  assign n2115 = n2114 ^ n1158;
  assign n2116 = n2115 ^ n1027;
  assign n2117 = n1881 & ~n2011;
  assign n2118 = n2117 ^ n1884;
  assign n2119 = n2118 ^ n2115;
  assign n2120 = n2116 & n2119;
  assign n2121 = n2120 ^ n1027;
  assign n2122 = n2121 ^ n905;
  assign n2123 = n1888 & ~n2011;
  assign n2124 = n2123 ^ n1890;
  assign n2125 = n2124 ^ n2121;
  assign n2126 = n2122 & ~n2125;
  assign n2127 = n2126 ^ n905;
  assign n2128 = n2127 ^ n803;
  assign n2129 = n1893 ^ n905;
  assign n2130 = ~n2011 & n2129;
  assign n2131 = n2130 ^ n1834;
  assign n2132 = n2131 ^ n2127;
  assign n2133 = n2128 & n2132;
  assign n2134 = n2133 ^ n803;
  assign n2135 = n2134 ^ n707;
  assign n2136 = n1896 ^ n803;
  assign n2137 = ~n2011 & n2136;
  assign n2138 = n2137 ^ n1830;
  assign n2139 = n2138 ^ n2134;
  assign n2140 = ~n2135 & ~n2139;
  assign n2141 = n2140 ^ n707;
  assign n2142 = n2141 ^ n608;
  assign n2143 = ~n1900 & ~n2011;
  assign n2144 = n2143 ^ n1906;
  assign n2145 = n2144 ^ n2141;
  assign n2146 = ~n2142 & ~n2145;
  assign n2147 = n2146 ^ n608;
  assign n2148 = n2147 ^ n514;
  assign n2149 = n1909 ^ n608;
  assign n2150 = ~n2011 & ~n2149;
  assign n2151 = n2150 ^ n1817;
  assign n2152 = n2151 ^ n2147;
  assign n2153 = n2148 & ~n2152;
  assign n2154 = n2153 ^ n514;
  assign n2155 = n2154 ^ n436;
  assign n2156 = n1909 ^ n1817;
  assign n2157 = ~n2149 & n2156;
  assign n2158 = n2157 ^ n608;
  assign n2159 = n2158 ^ n514;
  assign n2160 = ~n2011 & n2159;
  assign n2161 = n2160 ^ n1821;
  assign n2162 = n2161 ^ n2154;
  assign n2163 = n2155 & n2162;
  assign n2164 = n2163 ^ n436;
  assign n2165 = n2164 ^ n2052;
  assign n2166 = n2053 & ~n2165;
  assign n2167 = n2166 ^ n363;
  assign n2168 = n2167 ^ n2049;
  assign n2169 = ~n2050 & n2168;
  assign n2170 = n2169 ^ n300;
  assign n2171 = n2170 ^ n243;
  assign n2172 = n1938 & ~n2011;
  assign n2173 = n2172 ^ n1940;
  assign n2174 = n2173 ^ n2170;
  assign n2175 = n2171 & ~n2174;
  assign n2176 = n2175 ^ n243;
  assign n2177 = n2176 ^ n210;
  assign n2178 = n1944 & ~n2011;
  assign n2179 = n2178 ^ n1946;
  assign n2180 = n2179 ^ n2176;
  assign n2181 = n2177 & n2180;
  assign n2182 = n2181 ^ n210;
  assign n2183 = n2182 ^ n147;
  assign n2184 = n1950 & ~n2011;
  assign n2185 = n2184 ^ n1952;
  assign n2186 = n2185 ^ n2182;
  assign n2187 = ~n2183 & ~n2186;
  assign n2188 = n2187 ^ n147;
  assign n2189 = n2047 & n2188;
  assign n2190 = n132 & ~n2041;
  assign n2191 = ~n2038 & ~n2045;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = n2047 & ~n2192;
  assign n2194 = ~n2189 & ~n2193;
  assign n2195 = n2167 ^ n300;
  assign n2196 = n2194 & n2195;
  assign n2197 = n2196 ^ n2049;
  assign n2198 = n2197 ^ n243;
  assign n2199 = n2164 ^ n363;
  assign n2200 = n2194 & n2199;
  assign n2201 = n2200 ^ n2052;
  assign n2202 = n2201 ^ n300;
  assign n2203 = n2083 ^ n2011;
  assign n2204 = n2194 & ~n2203;
  assign n2205 = n2204 ^ n2011;
  assign n2206 = n2205 ^ x88;
  assign n2207 = n2206 ^ n1804;
  assign n2208 = ~x84 & ~x85;
  assign n2209 = ~n2011 & n2208;
  assign n2210 = ~x86 & n2209;
  assign n2211 = n2194 ^ x87;
  assign n2212 = n2011 & n2208;
  assign n2213 = ~x86 & n2212;
  assign n2214 = n2213 ^ n2011;
  assign n2215 = n2214 ^ n2194;
  assign n2216 = n2215 ^ n2214;
  assign n2217 = n2214 ^ x86;
  assign n2218 = n2217 ^ n2214;
  assign n2219 = n2216 & n2218;
  assign n2220 = n2219 ^ n2214;
  assign n2221 = n2211 & ~n2220;
  assign n2222 = n2221 ^ n2214;
  assign n2223 = ~n2210 & n2222;
  assign n2224 = n2223 ^ n2206;
  assign n2225 = ~n2207 & n2224;
  assign n2226 = n2225 ^ n1804;
  assign n2227 = n2226 ^ n1621;
  assign n2229 = n2087 ^ n2085;
  assign n2230 = n2229 ^ n2087;
  assign n2231 = n2089 ^ n2087;
  assign n2232 = n2231 ^ n2087;
  assign n2233 = ~n2230 & n2232;
  assign n2234 = n2233 ^ n2087;
  assign n2235 = n2011 & n2234;
  assign n2236 = n2235 ^ n2087;
  assign n2228 = ~x88 & ~n2011;
  assign n2237 = n2236 ^ n2228;
  assign n2238 = n2083 ^ n1804;
  assign n2239 = n2238 ^ n2236;
  assign n2240 = n2236 ^ n2194;
  assign n2241 = ~n2236 & ~n2240;
  assign n2242 = n2241 ^ n2236;
  assign n2243 = ~n2239 & ~n2242;
  assign n2244 = n2243 ^ n2241;
  assign n2245 = n2244 ^ n2236;
  assign n2246 = n2245 ^ n2194;
  assign n2247 = n2237 & ~n2246;
  assign n2248 = n2247 ^ n2228;
  assign n2249 = n2248 ^ x89;
  assign n2250 = n2249 ^ n2226;
  assign n2251 = n2227 & ~n2250;
  assign n2252 = n2251 ^ n1621;
  assign n2253 = n2252 ^ n1458;
  assign n2254 = n2099 & n2194;
  assign n2255 = n2254 ^ n2103;
  assign n2256 = n2255 ^ n2252;
  assign n2257 = n2253 & n2256;
  assign n2258 = n2257 ^ n1458;
  assign n2259 = n2258 ^ n1299;
  assign n2260 = n2106 ^ n1458;
  assign n2261 = n2194 & n2260;
  assign n2262 = n2261 ^ n2081;
  assign n2263 = n2262 ^ n2258;
  assign n2264 = n2259 & ~n2263;
  assign n2265 = n2264 ^ n1299;
  assign n2266 = n2265 ^ n1158;
  assign n2267 = n2109 ^ n1299;
  assign n2268 = n2194 & n2267;
  assign n2269 = n2268 ^ n2058;
  assign n2270 = n2269 ^ n2265;
  assign n2271 = n2266 & n2270;
  assign n2272 = n2271 ^ n1158;
  assign n2273 = n2272 ^ n1027;
  assign n2274 = n2112 ^ n1158;
  assign n2275 = n2194 & n2274;
  assign n2276 = n2275 ^ n2055;
  assign n2277 = n2276 ^ n2272;
  assign n2278 = n2273 & ~n2277;
  assign n2279 = n2278 ^ n1027;
  assign n2280 = n2279 ^ n905;
  assign n2281 = n2116 & n2194;
  assign n2282 = n2281 ^ n2118;
  assign n2283 = n2282 ^ n2279;
  assign n2284 = n2280 & n2283;
  assign n2285 = n2284 ^ n905;
  assign n2286 = n2285 ^ n803;
  assign n2287 = n2122 & n2194;
  assign n2288 = n2287 ^ n2124;
  assign n2289 = n2288 ^ n2285;
  assign n2290 = n2286 & ~n2289;
  assign n2291 = n2290 ^ n803;
  assign n2292 = n2291 ^ n707;
  assign n2293 = n2128 & n2194;
  assign n2294 = n2293 ^ n2131;
  assign n2295 = n2294 ^ n2291;
  assign n2296 = ~n2292 & n2295;
  assign n2297 = n2296 ^ n707;
  assign n2298 = n2297 ^ n608;
  assign n2299 = ~n2135 & n2194;
  assign n2300 = n2299 ^ n2138;
  assign n2301 = n2300 ^ n2297;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = n2302 ^ n608;
  assign n2304 = n2303 ^ n514;
  assign n2305 = ~n2142 & n2194;
  assign n2306 = n2305 ^ n2144;
  assign n2307 = n2306 ^ n2303;
  assign n2308 = n2304 & n2307;
  assign n2309 = n2308 ^ n514;
  assign n2310 = n2309 ^ n436;
  assign n2311 = n2148 & n2194;
  assign n2312 = n2311 ^ n2151;
  assign n2313 = n2312 ^ n2309;
  assign n2314 = n2310 & ~n2313;
  assign n2315 = n2314 ^ n436;
  assign n2316 = n2315 ^ n363;
  assign n2317 = n2155 & n2194;
  assign n2318 = n2317 ^ n2161;
  assign n2319 = n2318 ^ n2315;
  assign n2320 = n2316 & n2319;
  assign n2321 = n2320 ^ n363;
  assign n2322 = n2321 ^ n2201;
  assign n2323 = n2202 & ~n2322;
  assign n2324 = n2323 ^ n300;
  assign n2325 = n2324 ^ n2197;
  assign n2326 = ~n2198 & n2325;
  assign n2327 = n2326 ^ n243;
  assign n2328 = n2327 ^ n210;
  assign n2329 = n2171 & n2194;
  assign n2330 = n2329 ^ n2173;
  assign n2331 = n2330 ^ n2327;
  assign n2332 = n2328 & ~n2331;
  assign n2333 = n2332 ^ n210;
  assign n2334 = n2333 ^ n147;
  assign n2335 = n2041 & ~n2188;
  assign n2336 = n132 & n2335;
  assign n2337 = n2194 & n2336;
  assign n2338 = n133 & ~n2337;
  assign n2339 = ~n132 & ~n2189;
  assign n2340 = n2188 ^ n2041;
  assign n2341 = n2339 & ~n2340;
  assign n2342 = n2338 & ~n2341;
  assign n2343 = n2188 ^ n132;
  assign n2344 = n2041 ^ n132;
  assign n2345 = n2343 & ~n2344;
  assign n2346 = n2345 ^ n132;
  assign n2347 = ~n133 & ~n2346;
  assign n2348 = n2194 & n2347;
  assign n2349 = ~n2342 & ~n2348;
  assign n2350 = ~n2041 & ~n2194;
  assign n2351 = ~n2045 & ~n2350;
  assign n2352 = ~n2349 & n2351;
  assign n2353 = n2045 & ~n2348;
  assign n2354 = ~n2041 & n2188;
  assign n2355 = n1292 & n2354;
  assign n2356 = n2194 & n2355;
  assign n2357 = n2353 & ~n2356;
  assign n2358 = ~n2352 & ~n2357;
  assign n2359 = n2194 & n2343;
  assign n2360 = n2359 ^ n2041;
  assign n2361 = ~n133 & ~n2360;
  assign n2362 = n2177 & n2194;
  assign n2363 = n2362 ^ n2179;
  assign n2364 = n2363 ^ n2333;
  assign n2365 = ~n2334 & n2364;
  assign n2366 = n2365 ^ n147;
  assign n2367 = n2366 ^ n132;
  assign n2368 = ~n2183 & n2194;
  assign n2369 = n2368 ^ n2185;
  assign n2370 = n2369 ^ n2366;
  assign n2371 = n2367 & ~n2370;
  assign n2372 = n2371 ^ n2366;
  assign n2373 = ~n2361 & ~n2372;
  assign n2374 = n2358 & ~n2373;
  assign n2375 = ~n2334 & ~n2374;
  assign n2376 = n2375 ^ n2363;
  assign n2377 = n132 & n2376;
  assign n2378 = n2321 ^ n300;
  assign n2379 = ~n2374 & n2378;
  assign n2380 = n2379 ^ n2201;
  assign n2381 = n2380 ^ n243;
  assign n2382 = n2316 & ~n2374;
  assign n2383 = n2382 ^ n2318;
  assign n2384 = n2383 ^ n300;
  assign n2385 = n2266 & ~n2374;
  assign n2386 = n2385 ^ n2269;
  assign n2387 = n2386 ^ n1027;
  assign n2388 = n2259 & ~n2374;
  assign n2389 = n2388 ^ n2262;
  assign n2390 = n2389 ^ n1158;
  assign n2391 = n2227 & ~n2374;
  assign n2392 = n2391 ^ n2249;
  assign n2393 = n2392 ^ n1458;
  assign n2394 = n2223 ^ n1804;
  assign n2395 = ~n2374 & n2394;
  assign n2396 = n2395 ^ n2206;
  assign n2397 = n2396 ^ n1621;
  assign n2399 = n2194 ^ n2011;
  assign n2400 = n2399 ^ n2194;
  assign n2401 = n2400 ^ n2399;
  assign n2402 = n2399 ^ n2208;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = n2403 ^ n2399;
  assign n2405 = ~x86 & ~n2404;
  assign n2406 = n2405 ^ n2399;
  assign n2398 = ~x86 & n2194;
  assign n2407 = n2406 ^ n2398;
  assign n2408 = n2208 ^ n2011;
  assign n2409 = n2408 ^ n2406;
  assign n2410 = n2406 ^ n2374;
  assign n2411 = n2406 & ~n2410;
  assign n2412 = n2411 ^ n2406;
  assign n2413 = n2409 & n2412;
  assign n2414 = n2413 ^ n2411;
  assign n2415 = n2414 ^ n2406;
  assign n2416 = n2415 ^ n2374;
  assign n2417 = ~n2407 & ~n2416;
  assign n2418 = n2417 ^ n2398;
  assign n2419 = n2418 ^ x87;
  assign n2420 = n1804 & n2419;
  assign n2421 = n2420 ^ n2396;
  assign n2422 = ~n2397 & ~n2421;
  assign n2423 = n2422 ^ n2396;
  assign n2424 = n2423 ^ n2392;
  assign n2425 = n2424 ^ n2392;
  assign n2426 = ~n1804 & ~n2419;
  assign n2427 = ~n1621 & n2396;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = x84 & ~n2194;
  assign n2430 = ~x82 & ~x83;
  assign n2431 = ~n2194 & ~n2430;
  assign n2432 = ~n2429 & ~n2431;
  assign n2433 = n2374 ^ x85;
  assign n2434 = n2432 & n2433;
  assign n2436 = ~x85 & ~n2374;
  assign n2435 = n2194 & n2430;
  assign n2437 = n2436 ^ n2435;
  assign n2438 = x84 & n2437;
  assign n2439 = n2438 ^ n2435;
  assign n2440 = ~n2434 & ~n2439;
  assign n2441 = n2440 ^ n2011;
  assign n2442 = n2208 ^ n2194;
  assign n2443 = ~n2374 & n2442;
  assign n2444 = n2443 ^ n2194;
  assign n2445 = n2444 ^ x86;
  assign n2446 = n2445 ^ n2440;
  assign n2447 = n2441 & ~n2446;
  assign n2448 = n2447 ^ n2011;
  assign n2449 = n2428 & n2448;
  assign n2450 = n2449 ^ n2392;
  assign n2451 = n2450 ^ n2392;
  assign n2452 = n2425 & ~n2451;
  assign n2453 = n2452 ^ n2392;
  assign n2454 = n2393 & n2453;
  assign n2455 = n2454 ^ n1458;
  assign n2456 = n2455 ^ n1299;
  assign n2457 = n2253 & ~n2374;
  assign n2458 = n2457 ^ n2255;
  assign n2459 = n2458 ^ n2455;
  assign n2460 = n2456 & n2459;
  assign n2461 = n2460 ^ n1299;
  assign n2462 = n2461 ^ n2389;
  assign n2463 = n2390 & ~n2462;
  assign n2464 = n2463 ^ n1158;
  assign n2465 = n2464 ^ n2386;
  assign n2466 = ~n2387 & n2465;
  assign n2467 = n2466 ^ n1027;
  assign n2468 = n2467 ^ n905;
  assign n2469 = n2273 & ~n2374;
  assign n2470 = n2469 ^ n2276;
  assign n2471 = n2470 ^ n2467;
  assign n2472 = n2468 & ~n2471;
  assign n2473 = n2472 ^ n905;
  assign n2474 = n2473 ^ n803;
  assign n2475 = n2280 & ~n2374;
  assign n2476 = n2475 ^ n2282;
  assign n2477 = n2476 ^ n2473;
  assign n2478 = n2474 & n2477;
  assign n2479 = n2478 ^ n803;
  assign n2480 = n2479 ^ n707;
  assign n2481 = n2286 & ~n2374;
  assign n2482 = n2481 ^ n2288;
  assign n2483 = n2482 ^ n2479;
  assign n2484 = ~n2480 & ~n2483;
  assign n2485 = n2484 ^ n707;
  assign n2486 = n2485 ^ n608;
  assign n2487 = ~n2292 & ~n2374;
  assign n2488 = n2487 ^ n2294;
  assign n2489 = n2488 ^ n2485;
  assign n2490 = ~n2486 & ~n2489;
  assign n2491 = n2490 ^ n608;
  assign n2492 = n2491 ^ n514;
  assign n2493 = ~n2298 & ~n2374;
  assign n2494 = n2493 ^ n2300;
  assign n2495 = n2494 ^ n2491;
  assign n2496 = n2492 & ~n2495;
  assign n2497 = n2496 ^ n514;
  assign n2498 = n2497 ^ n436;
  assign n2499 = n2304 & ~n2374;
  assign n2500 = n2499 ^ n2306;
  assign n2501 = n2500 ^ n2497;
  assign n2502 = n2498 & n2501;
  assign n2503 = n2502 ^ n436;
  assign n2504 = n2503 ^ n363;
  assign n2505 = n2310 & ~n2374;
  assign n2506 = n2505 ^ n2312;
  assign n2507 = n2506 ^ n2503;
  assign n2508 = n2504 & ~n2507;
  assign n2509 = n2508 ^ n363;
  assign n2510 = n2509 ^ n2383;
  assign n2511 = ~n2384 & n2510;
  assign n2512 = n2511 ^ n300;
  assign n2513 = n2512 ^ n2380;
  assign n2514 = n2381 & ~n2513;
  assign n2515 = n2514 ^ n243;
  assign n2516 = n2515 ^ n210;
  assign n2517 = n2324 ^ n243;
  assign n2518 = ~n2374 & n2517;
  assign n2519 = n2518 ^ n2197;
  assign n2520 = n2519 ^ n2515;
  assign n2521 = n2516 & n2520;
  assign n2522 = n2521 ^ n210;
  assign n2523 = n2522 ^ n147;
  assign n2524 = n2328 & ~n2374;
  assign n2525 = n2524 ^ n2330;
  assign n2526 = n2525 ^ n2522;
  assign n2527 = ~n2523 & ~n2526;
  assign n2528 = n2527 ^ n147;
  assign n2529 = ~n2377 & ~n2528;
  assign n2530 = ~n132 & ~n2376;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = n132 & n2366;
  assign n2533 = ~n132 & ~n2366;
  assign n2534 = ~n2374 & ~n2533;
  assign n2535 = ~n2532 & n2534;
  assign n2536 = n2535 ^ n2369;
  assign n2537 = ~n2531 & n2536;
  assign n2561 = n2360 ^ n2358;
  assign n2562 = ~n2369 & ~n2533;
  assign n2563 = n2562 ^ n2358;
  assign n2564 = n2358 & ~n2563;
  assign n2565 = n2564 ^ n2358;
  assign n2566 = ~n2561 & n2565;
  assign n2567 = n2566 ^ n2564;
  assign n2568 = n2567 ^ n2358;
  assign n2569 = n2568 ^ n2562;
  assign n2570 = ~n2532 & ~n2569;
  assign n2571 = n2570 ^ n2360;
  assign n2538 = n2530 ^ n2360;
  assign n2539 = n2530 ^ n2372;
  assign n2540 = n2538 & n2539;
  assign n2541 = n2540 ^ n2371;
  assign n2542 = n2541 ^ n2366;
  assign n2543 = n2542 ^ n2360;
  assign n2544 = ~n2530 & n2543;
  assign n2545 = n2544 ^ n2530;
  assign n2546 = n2545 ^ n2369;
  assign n2547 = n2363 & n2366;
  assign n2548 = n2374 & n2547;
  assign n2549 = n2360 & n2532;
  assign n2550 = n132 & n2358;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2548 & n2551;
  assign n2553 = n2552 ^ n2545;
  assign n2554 = n2553 ^ n2552;
  assign n2555 = n2552 ^ n2534;
  assign n2556 = ~n2554 & n2555;
  assign n2557 = n2556 ^ n2552;
  assign n2558 = n2546 & n2557;
  assign n2559 = n2558 ^ n2369;
  assign n2560 = ~n2529 & ~n2559;
  assign n2572 = n2571 ^ n2560;
  assign n2573 = n2571 ^ n2358;
  assign n2574 = n2571 ^ n133;
  assign n2575 = n2571 & n2574;
  assign n2576 = n2575 ^ n2571;
  assign n2577 = n2573 & n2576;
  assign n2578 = n2577 ^ n2575;
  assign n2579 = n2578 ^ n2571;
  assign n2580 = n2579 ^ n133;
  assign n2581 = ~n2572 & n2580;
  assign n2582 = n2581 ^ n2571;
  assign n2583 = ~n2537 & ~n2582;
  assign n2584 = n2528 ^ n132;
  assign n2585 = ~n2583 & n2584;
  assign n2586 = n2585 ^ n2376;
  assign n2587 = ~n2523 & ~n2583;
  assign n2588 = n2587 ^ n2525;
  assign n2589 = n2516 & ~n2583;
  assign n2590 = n2589 ^ n2519;
  assign n2591 = n2590 ^ n147;
  assign n2592 = n2512 ^ n243;
  assign n2593 = ~n2583 & n2592;
  assign n2594 = n2593 ^ n2380;
  assign n2595 = n2594 ^ n210;
  assign n2596 = n2430 ^ n2374;
  assign n2597 = ~n2583 & ~n2596;
  assign n2598 = n2597 ^ n2374;
  assign n2599 = n2598 ^ x84;
  assign n2600 = n2599 ^ n2194;
  assign n2601 = ~x80 & ~x81;
  assign n2602 = ~n2374 & n2601;
  assign n2603 = ~x82 & n2602;
  assign n2604 = ~n2430 & ~n2583;
  assign n2605 = n2604 ^ x83;
  assign n2606 = n2604 ^ n2583;
  assign n2607 = n2374 & n2601;
  assign n2608 = ~x82 & n2607;
  assign n2609 = n2608 ^ n2374;
  assign n2610 = n2609 ^ n2583;
  assign n2611 = n2610 ^ n2583;
  assign n2612 = n2606 & n2611;
  assign n2613 = n2612 ^ n2583;
  assign n2614 = ~n2605 & ~n2613;
  assign n2615 = n2614 ^ x83;
  assign n2616 = ~n2603 & n2615;
  assign n2617 = n2616 ^ n2599;
  assign n2618 = n2600 & n2617;
  assign n2619 = n2618 ^ n2194;
  assign n2620 = n2619 ^ n2011;
  assign n2622 = ~x84 & n2430;
  assign n2623 = n2622 ^ n2194;
  assign n2624 = n2623 ^ n2429;
  assign n2625 = n2374 & n2624;
  assign n2626 = n2625 ^ n2429;
  assign n2621 = ~x84 & ~n2374;
  assign n2627 = n2626 ^ n2621;
  assign n2628 = n2430 ^ n2194;
  assign n2629 = n2628 ^ n2626;
  assign n2630 = n2626 ^ n2583;
  assign n2631 = ~n2626 & n2630;
  assign n2632 = n2631 ^ n2626;
  assign n2633 = n2629 & ~n2632;
  assign n2634 = n2633 ^ n2631;
  assign n2635 = n2634 ^ n2626;
  assign n2636 = n2635 ^ n2583;
  assign n2637 = n2627 & n2636;
  assign n2638 = n2637 ^ n2621;
  assign n2639 = n2638 ^ x85;
  assign n2640 = n2639 ^ n2619;
  assign n2641 = ~n2620 & n2640;
  assign n2642 = n2641 ^ n2011;
  assign n2643 = n2642 ^ n1804;
  assign n2644 = n2441 & ~n2583;
  assign n2645 = n2644 ^ n2445;
  assign n2646 = n2645 ^ n2642;
  assign n2647 = n2643 & ~n2646;
  assign n2648 = n2647 ^ n1804;
  assign n2649 = n2648 ^ n1621;
  assign n2650 = n2448 ^ n1804;
  assign n2651 = ~n2583 & n2650;
  assign n2652 = n2651 ^ n2419;
  assign n2653 = n2652 ^ n2648;
  assign n2654 = n2649 & ~n2653;
  assign n2655 = n2654 ^ n1621;
  assign n2656 = n2655 ^ n1458;
  assign n2657 = n2419 ^ n1804;
  assign n2658 = n2448 ^ n2419;
  assign n2659 = n2657 & ~n2658;
  assign n2660 = n2659 ^ n1804;
  assign n2661 = n2660 ^ n1621;
  assign n2662 = ~n2583 & n2661;
  assign n2663 = n2662 ^ n2396;
  assign n2664 = n2663 ^ n2655;
  assign n2665 = n2656 & n2664;
  assign n2666 = n2665 ^ n1458;
  assign n2667 = n2666 ^ n1299;
  assign n2668 = n2660 ^ n2396;
  assign n2669 = ~n2397 & n2668;
  assign n2670 = n2669 ^ n1621;
  assign n2671 = n2670 ^ n1458;
  assign n2672 = ~n2583 & n2671;
  assign n2673 = n2672 ^ n2392;
  assign n2674 = n2673 ^ n2666;
  assign n2675 = n2667 & ~n2674;
  assign n2676 = n2675 ^ n1299;
  assign n2677 = n2676 ^ n1158;
  assign n2678 = n2456 & ~n2583;
  assign n2679 = n2678 ^ n2458;
  assign n2680 = n2679 ^ n2676;
  assign n2681 = n2677 & n2680;
  assign n2682 = n2681 ^ n1158;
  assign n2683 = n2682 ^ n1027;
  assign n2684 = n2461 ^ n1158;
  assign n2685 = ~n2583 & n2684;
  assign n2686 = n2685 ^ n2389;
  assign n2687 = n2686 ^ n2682;
  assign n2688 = n2683 & ~n2687;
  assign n2689 = n2688 ^ n1027;
  assign n2690 = n2689 ^ n905;
  assign n2691 = n2464 ^ n1027;
  assign n2692 = ~n2583 & n2691;
  assign n2693 = n2692 ^ n2386;
  assign n2694 = n2693 ^ n2689;
  assign n2695 = n2690 & n2694;
  assign n2696 = n2695 ^ n905;
  assign n2697 = n2696 ^ n803;
  assign n2698 = n2468 & ~n2583;
  assign n2699 = n2698 ^ n2470;
  assign n2700 = n2699 ^ n2696;
  assign n2701 = n2697 & ~n2700;
  assign n2702 = n2701 ^ n803;
  assign n2703 = n2702 ^ n707;
  assign n2704 = n2474 & ~n2583;
  assign n2705 = n2704 ^ n2476;
  assign n2706 = n2705 ^ n2702;
  assign n2707 = ~n2703 & n2706;
  assign n2708 = n2707 ^ n707;
  assign n2709 = n2708 ^ n608;
  assign n2710 = ~n2480 & ~n2583;
  assign n2711 = n2710 ^ n2482;
  assign n2712 = n2711 ^ n2708;
  assign n2713 = ~n2709 & n2712;
  assign n2714 = n2713 ^ n608;
  assign n2715 = n2714 ^ n514;
  assign n2716 = ~n2486 & ~n2583;
  assign n2717 = n2716 ^ n2488;
  assign n2718 = n2717 ^ n2714;
  assign n2719 = n2715 & n2718;
  assign n2720 = n2719 ^ n514;
  assign n2721 = n2720 ^ n436;
  assign n2722 = n2492 & ~n2583;
  assign n2723 = n2722 ^ n2494;
  assign n2724 = n2723 ^ n2720;
  assign n2725 = n2721 & ~n2724;
  assign n2726 = n2725 ^ n436;
  assign n2727 = n2726 ^ n363;
  assign n2728 = n2498 & ~n2583;
  assign n2729 = n2728 ^ n2500;
  assign n2730 = n2729 ^ n2726;
  assign n2731 = n2727 & n2730;
  assign n2732 = n2731 ^ n363;
  assign n2733 = n2732 ^ n300;
  assign n2734 = n2504 & ~n2583;
  assign n2735 = n2734 ^ n2506;
  assign n2736 = n2735 ^ n2732;
  assign n2737 = n2733 & ~n2736;
  assign n2738 = n2737 ^ n300;
  assign n2739 = n2738 ^ n243;
  assign n2740 = n2509 ^ n300;
  assign n2741 = ~n2583 & n2740;
  assign n2742 = n2741 ^ n2383;
  assign n2743 = n2742 ^ n2738;
  assign n2744 = n2739 & n2743;
  assign n2745 = n2744 ^ n243;
  assign n2746 = n2745 ^ n2594;
  assign n2747 = n2595 & ~n2746;
  assign n2748 = n2747 ^ n210;
  assign n2749 = n2748 ^ n2590;
  assign n2750 = n2591 & n2749;
  assign n2751 = n2750 ^ n147;
  assign n2784 = ~n132 & ~n2751;
  assign n2752 = n2751 ^ n132;
  assign n2753 = ~n133 & n2586;
  assign n2754 = n2751 ^ n2588;
  assign n2755 = n2752 & n2754;
  assign n2756 = n2755 ^ n132;
  assign n2757 = ~n2753 & ~n2756;
  assign n2758 = n2376 & ~n2536;
  assign n2761 = ~n2536 & ~n2560;
  assign n2762 = n2584 & n2761;
  assign n2763 = n2377 & n2559;
  assign n2764 = n2528 & n2763;
  assign n2765 = ~n2762 & ~n2764;
  assign n2759 = n1287 & ~n2528;
  assign n2760 = n2582 & ~n2759;
  assign n2766 = n2765 ^ n2760;
  assign n2767 = n2766 ^ n2760;
  assign n2768 = n2760 ^ n133;
  assign n2769 = n2768 ^ n2760;
  assign n2770 = ~n2767 & n2769;
  assign n2771 = n2770 ^ n2760;
  assign n2772 = ~n2758 & ~n2771;
  assign n2773 = n2772 ^ n2760;
  assign n2774 = n133 & n2773;
  assign n2775 = ~n2531 & n2582;
  assign n2776 = n2529 & n2758;
  assign n2777 = n2776 ^ n2536;
  assign n2778 = ~n2775 & ~n2777;
  assign n2779 = ~n2537 & ~n2778;
  assign n2780 = n2773 & n2779;
  assign n2781 = ~n2774 & ~n2780;
  assign n2782 = ~n2757 & n2781;
  assign n2783 = n2752 & ~n2782;
  assign n2785 = n2784 ^ n2783;
  assign n2786 = ~n2588 & n2785;
  assign n2787 = n2786 ^ n2783;
  assign n2788 = n2586 & n2787;
  assign n2789 = ~n2588 & n2751;
  assign n2790 = n2782 & n2789;
  assign n2791 = ~n2788 & ~n2790;
  assign n2792 = n2739 & ~n2782;
  assign n2793 = n2792 ^ n2742;
  assign n2794 = n2793 ^ n210;
  assign n2795 = n2733 & ~n2782;
  assign n2796 = n2795 ^ n2735;
  assign n2797 = n2796 ^ n243;
  assign n2798 = n2616 ^ n2194;
  assign n2799 = ~n2782 & ~n2798;
  assign n2800 = n2799 ^ n2599;
  assign n2801 = n2800 ^ n2011;
  assign n2803 = n2583 ^ n2374;
  assign n2804 = n2803 ^ n2583;
  assign n2805 = n2804 ^ n2803;
  assign n2806 = n2803 ^ n2601;
  assign n2807 = n2805 & n2806;
  assign n2808 = n2807 ^ n2803;
  assign n2809 = ~x82 & n2808;
  assign n2810 = n2809 ^ n2803;
  assign n2802 = ~x82 & ~n2583;
  assign n2811 = n2810 ^ n2802;
  assign n2812 = n2601 ^ n2374;
  assign n2813 = n2812 ^ n2810;
  assign n2814 = n2810 ^ n2782;
  assign n2815 = ~n2810 & n2814;
  assign n2816 = n2815 ^ n2810;
  assign n2817 = ~n2813 & ~n2816;
  assign n2818 = n2817 ^ n2815;
  assign n2819 = n2818 ^ n2810;
  assign n2820 = n2819 ^ n2782;
  assign n2821 = n2811 & n2820;
  assign n2822 = n2821 ^ n2802;
  assign n2823 = n2822 ^ x83;
  assign n2824 = n2823 ^ n2194;
  assign n2825 = n2601 ^ n2583;
  assign n2826 = ~n2782 & ~n2825;
  assign n2827 = n2826 ^ n2583;
  assign n2828 = n2827 ^ x82;
  assign n2829 = n2828 ^ n2374;
  assign n2830 = n2782 ^ x81;
  assign n2831 = x80 & n2583;
  assign n2832 = ~x78 & ~x79;
  assign n2833 = n2583 & ~n2832;
  assign n2834 = ~n2831 & ~n2833;
  assign n2835 = n2830 & n2834;
  assign n2836 = ~n2583 & n2832;
  assign n2837 = n2836 ^ x81;
  assign n2838 = n2837 ^ n2836;
  assign n2839 = n2836 ^ n2782;
  assign n2840 = n2839 ^ n2836;
  assign n2841 = ~n2838 & ~n2840;
  assign n2842 = n2841 ^ n2836;
  assign n2843 = x80 & n2842;
  assign n2844 = n2843 ^ n2836;
  assign n2845 = ~n2835 & ~n2844;
  assign n2846 = n2845 ^ n2828;
  assign n2847 = ~n2829 & n2846;
  assign n2848 = n2847 ^ n2374;
  assign n2849 = n2848 ^ n2823;
  assign n2850 = ~n2824 & ~n2849;
  assign n2851 = n2850 ^ n2194;
  assign n2852 = n2851 ^ n2800;
  assign n2853 = ~n2801 & ~n2852;
  assign n2854 = n2853 ^ n2011;
  assign n2855 = n2854 ^ n1804;
  assign n2856 = ~n2620 & ~n2782;
  assign n2857 = n2856 ^ n2639;
  assign n2858 = n2857 ^ n2854;
  assign n2859 = n2855 & ~n2858;
  assign n2860 = n2859 ^ n1804;
  assign n2861 = n2860 ^ n1621;
  assign n2862 = n2643 & ~n2782;
  assign n2863 = n2862 ^ n2645;
  assign n2864 = n2863 ^ n2860;
  assign n2865 = n2861 & ~n2864;
  assign n2866 = n2865 ^ n1621;
  assign n2867 = n2866 ^ n1458;
  assign n2868 = n2649 & ~n2782;
  assign n2869 = n2868 ^ n2652;
  assign n2870 = n2869 ^ n2866;
  assign n2871 = n2867 & ~n2870;
  assign n2872 = n2871 ^ n1458;
  assign n2873 = n2872 ^ n1299;
  assign n2874 = n2656 & ~n2782;
  assign n2875 = n2874 ^ n2663;
  assign n2876 = n2875 ^ n2872;
  assign n2877 = n2873 & n2876;
  assign n2878 = n2877 ^ n1299;
  assign n2879 = n2878 ^ n1158;
  assign n2880 = n2667 & ~n2782;
  assign n2881 = n2880 ^ n2673;
  assign n2882 = n2881 ^ n2878;
  assign n2883 = n2879 & ~n2882;
  assign n2884 = n2883 ^ n1158;
  assign n2885 = n2884 ^ n1027;
  assign n2886 = n2677 & ~n2782;
  assign n2887 = n2886 ^ n2679;
  assign n2888 = n2887 ^ n2884;
  assign n2889 = n2885 & n2888;
  assign n2890 = n2889 ^ n1027;
  assign n2891 = n2890 ^ n905;
  assign n2892 = n2683 & ~n2782;
  assign n2893 = n2892 ^ n2686;
  assign n2894 = n2893 ^ n2890;
  assign n2895 = n2891 & ~n2894;
  assign n2896 = n2895 ^ n905;
  assign n2897 = n2896 ^ n803;
  assign n2898 = n2690 & ~n2782;
  assign n2899 = n2898 ^ n2693;
  assign n2900 = n2899 ^ n2896;
  assign n2901 = n2897 & n2900;
  assign n2902 = n2901 ^ n803;
  assign n2903 = n2902 ^ n707;
  assign n2904 = n2697 & ~n2782;
  assign n2905 = n2904 ^ n2699;
  assign n2906 = n2905 ^ n2902;
  assign n2907 = ~n2903 & ~n2906;
  assign n2908 = n2907 ^ n707;
  assign n2909 = n2908 ^ n608;
  assign n2910 = ~n2703 & ~n2782;
  assign n2911 = n2910 ^ n2705;
  assign n2912 = n2911 ^ n2908;
  assign n2913 = ~n2909 & ~n2912;
  assign n2914 = n2913 ^ n608;
  assign n2915 = n2914 ^ n514;
  assign n2916 = ~n2709 & ~n2782;
  assign n2917 = n2916 ^ n2711;
  assign n2918 = n2917 ^ n2914;
  assign n2919 = n2915 & ~n2918;
  assign n2920 = n2919 ^ n514;
  assign n2921 = n2920 ^ n436;
  assign n2922 = n2715 & ~n2782;
  assign n2923 = n2922 ^ n2717;
  assign n2924 = n2923 ^ n2920;
  assign n2925 = n2921 & n2924;
  assign n2926 = n2925 ^ n436;
  assign n2927 = n2926 ^ n363;
  assign n2928 = n2721 & ~n2782;
  assign n2929 = n2928 ^ n2723;
  assign n2930 = n2929 ^ n2926;
  assign n2931 = n2927 & ~n2930;
  assign n2932 = n2931 ^ n363;
  assign n2933 = n2932 ^ n300;
  assign n2934 = n2727 & ~n2782;
  assign n2935 = n2934 ^ n2729;
  assign n2936 = n2935 ^ n2932;
  assign n2937 = n2933 & n2936;
  assign n2938 = n2937 ^ n300;
  assign n2939 = n2938 ^ n2796;
  assign n2940 = n2797 & ~n2939;
  assign n2941 = n2940 ^ n243;
  assign n2942 = n2941 ^ n2793;
  assign n2943 = ~n2794 & n2942;
  assign n2944 = n2943 ^ n210;
  assign n2945 = n2944 ^ n147;
  assign n2946 = n2745 ^ n210;
  assign n2947 = ~n2782 & n2946;
  assign n2948 = n2947 ^ n2594;
  assign n2949 = n2948 ^ n2944;
  assign n2950 = ~n2945 & ~n2949;
  assign n2951 = n2950 ^ n147;
  assign n2952 = ~n2791 & n2951;
  assign n2953 = n2588 ^ n2586;
  assign n2954 = n2754 & ~n2953;
  assign n2955 = n2954 ^ n2588;
  assign n2956 = ~n2782 & ~n2955;
  assign n2957 = n2956 ^ n2588;
  assign n2958 = n132 & ~n2957;
  assign n2959 = ~n2952 & ~n2958;
  assign n2960 = n2748 ^ n147;
  assign n2961 = ~n2782 & ~n2960;
  assign n2962 = n2961 ^ n2590;
  assign n2963 = ~n2951 & ~n2962;
  assign n2964 = ~n132 & ~n2962;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = ~n2959 & n2965;
  assign n2967 = n133 & ~n2966;
  assign n2969 = n2753 & n2780;
  assign n2968 = ~n2586 & ~n2774;
  assign n2970 = n2969 ^ n2968;
  assign n2971 = ~n2756 & n2970;
  assign n2972 = n2971 ^ n2968;
  assign n2973 = ~n2967 & ~n2972;
  assign n2974 = n2783 ^ n2588;
  assign n2975 = n2951 ^ n132;
  assign n2976 = n2962 ^ n2951;
  assign n2977 = n2975 & ~n2976;
  assign n2978 = n2977 ^ n132;
  assign n2979 = n2974 & ~n2978;
  assign n2980 = n2973 & ~n2979;
  assign n2981 = n2980 ^ x79;
  assign n2982 = ~x76 & ~x77;
  assign n2983 = n2782 & n2982;
  assign n2984 = ~x78 & n2983;
  assign n2985 = n2984 ^ n2782;
  assign n2986 = n2981 & ~n2985;
  assign n2987 = ~n2782 & n2982;
  assign n2988 = n2987 ^ x79;
  assign n2989 = n2988 ^ n2987;
  assign n2990 = n2987 ^ n2980;
  assign n2991 = n2990 ^ n2987;
  assign n2992 = ~n2989 & ~n2991;
  assign n2993 = n2992 ^ n2987;
  assign n2994 = x78 & n2993;
  assign n2995 = n2994 ^ n2987;
  assign n2996 = ~n2986 & ~n2995;
  assign n2997 = n2996 ^ n2583;
  assign n2998 = n2832 ^ n2782;
  assign n2999 = ~n2980 & ~n2998;
  assign n3000 = n2999 ^ n2782;
  assign n3001 = n3000 ^ x80;
  assign n3002 = n3001 ^ n2996;
  assign n3003 = n2997 & n3002;
  assign n3004 = n3003 ^ n2583;
  assign n3005 = n3004 ^ n2374;
  assign n3007 = ~x80 & n2832;
  assign n3008 = n3007 ^ n2583;
  assign n3009 = n3008 ^ n2831;
  assign n3010 = n2782 & ~n3009;
  assign n3011 = n3010 ^ n2831;
  assign n3006 = ~x80 & ~n2782;
  assign n3012 = n3011 ^ n3006;
  assign n3013 = n2832 ^ n2583;
  assign n3014 = n3013 ^ n3011;
  assign n3015 = n3011 ^ n2980;
  assign n3016 = ~n3011 & n3015;
  assign n3017 = n3016 ^ n3011;
  assign n3018 = ~n3014 & ~n3017;
  assign n3019 = n3018 ^ n3016;
  assign n3020 = n3019 ^ n3011;
  assign n3021 = n3020 ^ n2980;
  assign n3022 = n3012 & n3021;
  assign n3023 = n3022 ^ n3006;
  assign n3024 = n3023 ^ x81;
  assign n3025 = n3024 ^ n3004;
  assign n3026 = n3005 & ~n3025;
  assign n3027 = n3026 ^ n2374;
  assign n3028 = n3027 ^ n2194;
  assign n3029 = n2845 ^ n2374;
  assign n3030 = ~n2980 & n3029;
  assign n3031 = n3030 ^ n2828;
  assign n3032 = n3031 ^ n3027;
  assign n3033 = ~n3028 & n3032;
  assign n3034 = n3033 ^ n2194;
  assign n3035 = n3034 ^ n2011;
  assign n3036 = n2975 & ~n2980;
  assign n3037 = n3036 ^ n2962;
  assign n3038 = ~n133 & n3037;
  assign n3039 = n2897 & ~n2980;
  assign n3040 = n3039 ^ n2899;
  assign n3041 = n707 & n3040;
  assign n3042 = ~n2903 & ~n2980;
  assign n3043 = n3042 ^ n2905;
  assign n3044 = ~n608 & ~n3043;
  assign n3045 = ~n3041 & ~n3044;
  assign n3046 = n2861 & ~n2980;
  assign n3047 = n3046 ^ n2863;
  assign n3048 = n3047 ^ n1458;
  assign n3049 = n2855 & ~n2980;
  assign n3050 = n3049 ^ n2857;
  assign n3051 = n3050 ^ n1621;
  assign n3052 = n2848 ^ n2194;
  assign n3053 = ~n2980 & ~n3052;
  assign n3054 = n3053 ^ n2823;
  assign n3055 = n3054 ^ n3034;
  assign n3056 = ~n3035 & n3055;
  assign n3057 = n3056 ^ n2011;
  assign n3058 = n3057 ^ n1804;
  assign n3059 = n2851 ^ n2011;
  assign n3060 = ~n2980 & ~n3059;
  assign n3061 = n3060 ^ n2800;
  assign n3062 = n3061 ^ n3057;
  assign n3063 = n3058 & n3062;
  assign n3064 = n3063 ^ n1804;
  assign n3065 = n3064 ^ n3050;
  assign n3066 = n3051 & ~n3065;
  assign n3067 = n3066 ^ n1621;
  assign n3068 = n3067 ^ n3047;
  assign n3069 = n3048 & ~n3068;
  assign n3070 = n3069 ^ n1458;
  assign n3071 = n3070 ^ n1299;
  assign n3072 = n2867 & ~n2980;
  assign n3073 = n3072 ^ n2869;
  assign n3074 = n3073 ^ n3070;
  assign n3075 = n3071 & ~n3074;
  assign n3076 = n3075 ^ n1299;
  assign n3077 = n3076 ^ n1158;
  assign n3078 = n2873 & ~n2980;
  assign n3079 = n3078 ^ n2875;
  assign n3080 = n3079 ^ n3076;
  assign n3081 = n3077 & n3080;
  assign n3082 = n3081 ^ n1158;
  assign n3083 = n3082 ^ n1027;
  assign n3084 = n2879 & ~n2980;
  assign n3085 = n3084 ^ n2881;
  assign n3086 = n3085 ^ n3082;
  assign n3087 = n3083 & ~n3086;
  assign n3088 = n3087 ^ n1027;
  assign n3089 = n3088 ^ n905;
  assign n3090 = n2885 & ~n2980;
  assign n3091 = n3090 ^ n2887;
  assign n3092 = n3091 ^ n3088;
  assign n3093 = n3089 & n3092;
  assign n3094 = n3093 ^ n905;
  assign n3095 = n3094 ^ n803;
  assign n3096 = n2891 & ~n2980;
  assign n3097 = n3096 ^ n2893;
  assign n3098 = n3097 ^ n3094;
  assign n3099 = n3095 & ~n3098;
  assign n3100 = n3099 ^ n803;
  assign n3101 = n3045 & n3100;
  assign n3102 = n3043 ^ n608;
  assign n3103 = ~n707 & ~n3040;
  assign n3104 = n3103 ^ n3043;
  assign n3105 = n3102 & ~n3104;
  assign n3106 = n3105 ^ n608;
  assign n3107 = ~n3101 & ~n3106;
  assign n3108 = n3107 ^ n514;
  assign n3109 = ~n2909 & ~n2980;
  assign n3110 = n3109 ^ n2911;
  assign n3111 = n3110 ^ n3107;
  assign n3112 = ~n3108 & ~n3111;
  assign n3113 = n3112 ^ n514;
  assign n3114 = n3113 ^ n436;
  assign n3115 = n2915 & ~n2980;
  assign n3116 = n3115 ^ n2917;
  assign n3117 = n3116 ^ n3113;
  assign n3118 = n3114 & ~n3117;
  assign n3119 = n3118 ^ n436;
  assign n3120 = n3119 ^ n363;
  assign n3121 = n2921 & ~n2980;
  assign n3122 = n3121 ^ n2923;
  assign n3123 = n3122 ^ n3119;
  assign n3124 = n3120 & n3123;
  assign n3125 = n3124 ^ n363;
  assign n3126 = n3125 ^ n300;
  assign n3127 = n2927 & ~n2980;
  assign n3128 = n3127 ^ n2929;
  assign n3129 = n3128 ^ n3125;
  assign n3130 = n3126 & ~n3129;
  assign n3131 = n3130 ^ n300;
  assign n3132 = n3131 ^ n243;
  assign n3133 = n2933 & ~n2980;
  assign n3134 = n3133 ^ n2935;
  assign n3135 = n3134 ^ n3131;
  assign n3136 = n3132 & n3135;
  assign n3137 = n3136 ^ n243;
  assign n3138 = n3137 ^ n210;
  assign n3139 = n2938 ^ n243;
  assign n3140 = ~n2980 & n3139;
  assign n3141 = n3140 ^ n2796;
  assign n3142 = n3141 ^ n3137;
  assign n3143 = n3138 & ~n3142;
  assign n3144 = n3143 ^ n210;
  assign n3145 = n3144 ^ n147;
  assign n3146 = n2941 ^ n210;
  assign n3147 = ~n2980 & n3146;
  assign n3148 = n3147 ^ n2793;
  assign n3149 = n3148 ^ n3144;
  assign n3150 = ~n3145 & n3149;
  assign n3151 = n3150 ^ n147;
  assign n3152 = n3151 ^ n132;
  assign n3153 = ~n2945 & ~n2980;
  assign n3154 = n3153 ^ n2948;
  assign n3155 = n3154 ^ n3151;
  assign n3156 = n3152 & n3155;
  assign n3157 = n3156 ^ n132;
  assign n3158 = ~n3038 & ~n3157;
  assign n3159 = n2962 & n2980;
  assign n3160 = ~n2972 & ~n2974;
  assign n3161 = n3160 ^ n133;
  assign n3162 = n3161 ^ n3160;
  assign n3163 = ~n132 & n2963;
  assign n3164 = n3163 ^ n3160;
  assign n3165 = n3162 & n3164;
  assign n3166 = n3165 ^ n3160;
  assign n3167 = ~n2978 & ~n3166;
  assign n3168 = n3167 ^ n133;
  assign n3169 = ~n2974 & n3168;
  assign n3170 = ~n3159 & n3169;
  assign n3171 = ~n133 & ~n2978;
  assign n3172 = n2951 & n2962;
  assign n3173 = n1292 & n3172;
  assign n3174 = n2974 & ~n3173;
  assign n3175 = ~n3171 & n3174;
  assign n3176 = ~n3170 & ~n3175;
  assign n3177 = ~n3158 & n3176;
  assign n3178 = ~n3035 & ~n3177;
  assign n3179 = n3178 ^ n3054;
  assign n3180 = n3179 ^ n1804;
  assign n3181 = ~n3028 & ~n3177;
  assign n3182 = n3181 ^ n3031;
  assign n3183 = n3182 ^ n2011;
  assign n3184 = n3005 & ~n3177;
  assign n3185 = n3184 ^ n3024;
  assign n3186 = n3185 ^ n2194;
  assign n3245 = n2997 & ~n3177;
  assign n3246 = n3245 ^ n3001;
  assign n3187 = ~x74 & ~x75;
  assign n3191 = ~n2980 & n3187;
  assign n3192 = n2982 & ~n3191;
  assign n3188 = ~x76 & n3187;
  assign n3189 = x77 & ~n3188;
  assign n3190 = ~n2980 & n3189;
  assign n3193 = n3192 ^ n3190;
  assign n3194 = ~n3177 & n3193;
  assign n3195 = n3194 ^ n3190;
  assign n3196 = ~x78 & n3195;
  assign n3197 = ~n3177 & ~n3189;
  assign n3198 = ~x77 & n3188;
  assign n3199 = x78 & ~n3198;
  assign n3200 = n2980 & n3199;
  assign n3201 = ~n3197 & n3200;
  assign n3202 = ~n2782 & ~n3201;
  assign n3203 = ~n3196 & n3202;
  assign n3204 = x78 & ~n2980;
  assign n3205 = n3188 ^ x77;
  assign n3206 = n3177 ^ x77;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = n3207 ^ x77;
  assign n3209 = n3204 & ~n3208;
  assign n3210 = ~n3203 & ~n3209;
  assign n3211 = n2980 & n3177;
  assign n3212 = n3198 & n3211;
  assign n3213 = ~n2982 & ~n3177;
  assign n3214 = n2980 & n3189;
  assign n3215 = n3213 & ~n3214;
  assign n3216 = ~n3212 & ~n3215;
  assign n3217 = ~x78 & ~n3216;
  assign n3218 = n3210 & ~n3217;
  assign n3219 = n3218 ^ n2583;
  assign n3221 = n2980 ^ n2782;
  assign n3222 = n3221 ^ n2980;
  assign n3223 = n3222 ^ n3221;
  assign n3224 = n3221 ^ n2982;
  assign n3225 = n3223 & n3224;
  assign n3226 = n3225 ^ n3221;
  assign n3227 = ~x78 & n3226;
  assign n3228 = n3227 ^ n3221;
  assign n3220 = ~x78 & ~n2980;
  assign n3229 = n3228 ^ n3220;
  assign n3230 = n2982 ^ n2782;
  assign n3231 = n3230 ^ n3228;
  assign n3232 = n3228 ^ n3177;
  assign n3233 = ~n3228 & n3232;
  assign n3234 = n3233 ^ n3228;
  assign n3235 = ~n3231 & ~n3234;
  assign n3236 = n3235 ^ n3233;
  assign n3237 = n3236 ^ n3228;
  assign n3238 = n3237 ^ n3177;
  assign n3239 = n3229 & n3238;
  assign n3240 = n3239 ^ n3220;
  assign n3241 = n3240 ^ x79;
  assign n3242 = n3241 ^ n3218;
  assign n3243 = n3219 & ~n3242;
  assign n3244 = n3243 ^ n2583;
  assign n3247 = n3246 ^ n3244;
  assign n3248 = n3246 ^ n2374;
  assign n3249 = n3247 & ~n3248;
  assign n3250 = n3249 ^ n2374;
  assign n3251 = n3250 ^ n3185;
  assign n3252 = ~n3186 & ~n3251;
  assign n3253 = n3252 ^ n2194;
  assign n3254 = n3253 ^ n3182;
  assign n3255 = ~n3183 & ~n3254;
  assign n3256 = n3255 ^ n2011;
  assign n3257 = n3256 ^ n3179;
  assign n3258 = n3180 & ~n3257;
  assign n3259 = n3258 ^ n1804;
  assign n3260 = n3259 ^ n1621;
  assign n3261 = n3058 & ~n3177;
  assign n3262 = n3261 ^ n3061;
  assign n3263 = n3262 ^ n3259;
  assign n3264 = n3260 & n3263;
  assign n3265 = n3264 ^ n1621;
  assign n3266 = n3265 ^ n1458;
  assign n3267 = n3064 ^ n1621;
  assign n3268 = ~n3177 & n3267;
  assign n3269 = n3268 ^ n3050;
  assign n3270 = n3269 ^ n3265;
  assign n3271 = n3266 & ~n3270;
  assign n3272 = n3271 ^ n1458;
  assign n3273 = n3272 ^ n1299;
  assign n3274 = n3067 ^ n1458;
  assign n3275 = ~n3177 & n3274;
  assign n3276 = n3275 ^ n3047;
  assign n3277 = n3276 ^ n3272;
  assign n3278 = n3273 & ~n3277;
  assign n3279 = n3278 ^ n1299;
  assign n3280 = n3279 ^ n1158;
  assign n3281 = n3071 & ~n3177;
  assign n3282 = n3281 ^ n3073;
  assign n3283 = n3282 ^ n3279;
  assign n3284 = n3280 & ~n3283;
  assign n3285 = n3284 ^ n1158;
  assign n3286 = n3285 ^ n1027;
  assign n3287 = n3077 & ~n3177;
  assign n3288 = n3287 ^ n3079;
  assign n3289 = n3288 ^ n3285;
  assign n3290 = n3286 & n3289;
  assign n3291 = n3290 ^ n1027;
  assign n3292 = n3291 ^ n905;
  assign n3293 = n3083 & ~n3177;
  assign n3294 = n3293 ^ n3085;
  assign n3295 = n3294 ^ n3291;
  assign n3296 = n3292 & ~n3295;
  assign n3297 = n3296 ^ n905;
  assign n3298 = n3297 ^ n803;
  assign n3299 = n3089 & ~n3177;
  assign n3300 = n3299 ^ n3091;
  assign n3301 = n3300 ^ n3297;
  assign n3302 = n3298 & n3301;
  assign n3303 = n3302 ^ n803;
  assign n3304 = n3303 ^ n707;
  assign n3305 = n3095 & ~n3177;
  assign n3306 = n3305 ^ n3097;
  assign n3307 = n3306 ^ n3303;
  assign n3308 = ~n3304 & ~n3307;
  assign n3309 = n3308 ^ n707;
  assign n3310 = n3309 ^ n608;
  assign n3311 = n3100 ^ n707;
  assign n3312 = ~n3177 & ~n3311;
  assign n3313 = n3312 ^ n3040;
  assign n3314 = n3313 ^ n3309;
  assign n3315 = ~n3310 & ~n3314;
  assign n3316 = n3315 ^ n608;
  assign n3317 = n3316 ^ n514;
  assign n3318 = n3100 ^ n3040;
  assign n3319 = ~n3311 & n3318;
  assign n3320 = n3319 ^ n707;
  assign n3321 = n3320 ^ n608;
  assign n3322 = ~n3177 & ~n3321;
  assign n3323 = n3322 ^ n3043;
  assign n3324 = n3323 ^ n3316;
  assign n3325 = n3317 & ~n3324;
  assign n3326 = n3325 ^ n514;
  assign n3327 = n3326 ^ n436;
  assign n3328 = ~n3108 & ~n3177;
  assign n3329 = n3328 ^ n3110;
  assign n3330 = n3329 ^ n3326;
  assign n3331 = n3327 & n3330;
  assign n3332 = n3331 ^ n436;
  assign n3333 = n3332 ^ n363;
  assign n3334 = n3114 & ~n3177;
  assign n3335 = n3334 ^ n3116;
  assign n3336 = n3335 ^ n3332;
  assign n3337 = n3333 & ~n3336;
  assign n3338 = n3337 ^ n363;
  assign n3339 = n3338 ^ n300;
  assign n3340 = ~n3145 & ~n3177;
  assign n3341 = n3340 ^ n3148;
  assign n3342 = n3120 & ~n3177;
  assign n3343 = n3342 ^ n3122;
  assign n3344 = n3343 ^ n3338;
  assign n3345 = n3339 & n3344;
  assign n3346 = n3345 ^ n300;
  assign n3347 = n3346 ^ n243;
  assign n3348 = n3126 & ~n3177;
  assign n3349 = n3348 ^ n3128;
  assign n3350 = n3349 ^ n3346;
  assign n3351 = n3347 & ~n3350;
  assign n3352 = n3351 ^ n243;
  assign n3353 = n3352 ^ n210;
  assign n3354 = n3132 & ~n3177;
  assign n3355 = n3354 ^ n3134;
  assign n3356 = n3355 ^ n3352;
  assign n3357 = n3353 & n3356;
  assign n3358 = n3357 ^ n210;
  assign n3359 = n3358 ^ n147;
  assign n3360 = n3138 & ~n3177;
  assign n3361 = n3360 ^ n3141;
  assign n3362 = n3361 ^ n3358;
  assign n3363 = ~n3359 & ~n3362;
  assign n3364 = n3363 ^ n147;
  assign n3365 = ~n3341 & ~n3364;
  assign n3366 = n1292 & ~n3154;
  assign n3367 = n3151 & n3366;
  assign n3368 = ~n3365 & n3367;
  assign n3369 = ~n133 & ~n3157;
  assign n3370 = ~n3368 & ~n3369;
  assign n3371 = ~n3037 & ~n3177;
  assign n3372 = ~n3370 & n3371;
  assign n3373 = ~n3154 & n3176;
  assign n3374 = n3154 ^ n3152;
  assign n3375 = n3154 ^ n133;
  assign n3376 = ~n3154 & ~n3375;
  assign n3377 = n3376 ^ n3154;
  assign n3378 = ~n3155 & ~n3377;
  assign n3379 = n3378 ^ n3376;
  assign n3380 = n3379 ^ n3154;
  assign n3381 = n3380 ^ n133;
  assign n3382 = ~n3374 & ~n3381;
  assign n3383 = ~n3373 & ~n3382;
  assign n3384 = n3037 & ~n3383;
  assign n3385 = n3364 ^ n132;
  assign n3386 = n3364 ^ n3341;
  assign n3387 = n3385 & ~n3386;
  assign n3388 = n3387 ^ n132;
  assign n3389 = n3384 & n3388;
  assign n3390 = ~n3157 & ~n3176;
  assign n3391 = n3038 & ~n3390;
  assign n3392 = ~n3389 & ~n3391;
  assign n3393 = ~n3372 & n3392;
  assign n3394 = n3152 & ~n3177;
  assign n3395 = n3394 ^ n3154;
  assign n3396 = ~n3388 & n3395;
  assign n3397 = ~n3393 & ~n3396;
  assign n3398 = n3339 & ~n3397;
  assign n3399 = n3398 ^ n3343;
  assign n3400 = ~n243 & n3399;
  assign n3401 = n3347 & ~n3397;
  assign n3402 = n3401 ^ n3349;
  assign n3403 = ~n210 & ~n3402;
  assign n3404 = ~n3400 & ~n3403;
  assign n3405 = n3317 & ~n3397;
  assign n3406 = n3405 ^ n3323;
  assign n3407 = n3406 ^ n436;
  assign n3569 = ~n3310 & ~n3397;
  assign n3570 = n3569 ^ n3313;
  assign n3408 = n3292 & ~n3397;
  assign n3409 = n3408 ^ n3294;
  assign n3410 = n3409 ^ n803;
  assign n3411 = n3286 & ~n3397;
  assign n3412 = n3411 ^ n3288;
  assign n3413 = n3412 ^ n905;
  assign n3414 = n3250 ^ n2194;
  assign n3415 = ~n3397 & ~n3414;
  assign n3416 = n3415 ^ n3185;
  assign n3417 = n3416 ^ n2011;
  assign n3429 = ~n3211 & ~n3213;
  assign n3430 = n3429 ^ x78;
  assign n3418 = ~n2980 & n3188;
  assign n3419 = x76 & ~n3177;
  assign n3420 = ~x77 & n3419;
  assign n3421 = ~n3418 & ~n3420;
  assign n3422 = x76 & n2980;
  assign n3423 = n2980 & ~n3187;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = n3206 & n3424;
  assign n3426 = n3421 & ~n3425;
  assign n3427 = n3426 ^ n2782;
  assign n3428 = ~n3397 & n3427;
  assign n3431 = n3430 ^ n3428;
  assign n3432 = n3431 ^ n2583;
  assign n3433 = x75 & ~n3397;
  assign n3434 = n3177 & ~n3433;
  assign n3435 = ~x72 & ~x73;
  assign n3436 = ~x74 & n3435;
  assign n3437 = ~n3434 & n3436;
  assign n3438 = n3397 & ~n3436;
  assign n3439 = ~x75 & x76;
  assign n3440 = ~n3438 & n3439;
  assign n3441 = ~n3419 & ~n3440;
  assign n3442 = ~n3437 & n3441;
  assign n3443 = ~n3177 & n3397;
  assign n3444 = x75 & n3443;
  assign n3445 = n3187 & ~n3397;
  assign n3446 = ~x76 & ~n3445;
  assign n3447 = ~n3444 & n3446;
  assign n3448 = n3442 & ~n3447;
  assign n3449 = ~n3177 & n3436;
  assign n3450 = n3439 & n3449;
  assign n3451 = n2980 & ~n3450;
  assign n3452 = n3188 & n3435;
  assign n3453 = n3452 ^ x76;
  assign n3454 = n3453 ^ n3452;
  assign n3455 = x75 & ~n3436;
  assign n3456 = n3455 ^ n3452;
  assign n3457 = n3456 ^ n3452;
  assign n3458 = n3454 & ~n3457;
  assign n3459 = n3458 ^ n3452;
  assign n3460 = ~n3177 & n3459;
  assign n3461 = n3460 ^ n3452;
  assign n3462 = n3461 ^ n3397;
  assign n3463 = n3462 ^ n3461;
  assign n3464 = n3177 & n3455;
  assign n3465 = ~x76 & ~n3187;
  assign n3466 = ~n3464 & n3465;
  assign n3467 = n3466 ^ n3461;
  assign n3468 = ~n3463 & n3467;
  assign n3469 = n3468 ^ n3461;
  assign n3470 = n3451 & ~n3469;
  assign n3471 = ~n3448 & ~n3470;
  assign n3472 = n3471 ^ n2782;
  assign n3474 = ~n3418 & n3424;
  assign n3475 = n3474 ^ n3422;
  assign n3476 = n3177 & n3475;
  assign n3477 = n3476 ^ n3422;
  assign n3473 = ~x76 & ~n3177;
  assign n3478 = n3477 ^ n3473;
  assign n3479 = n3187 ^ n2980;
  assign n3480 = n3479 ^ n3477;
  assign n3481 = n3477 ^ n3397;
  assign n3482 = ~n3477 & n3481;
  assign n3483 = n3482 ^ n3477;
  assign n3484 = ~n3480 & ~n3483;
  assign n3485 = n3484 ^ n3482;
  assign n3486 = n3485 ^ n3477;
  assign n3487 = n3486 ^ n3397;
  assign n3488 = n3478 & n3487;
  assign n3489 = n3488 ^ n3473;
  assign n3490 = n3489 ^ x77;
  assign n3491 = n3490 ^ n3471;
  assign n3492 = ~n3472 & n3491;
  assign n3493 = n3492 ^ n2782;
  assign n3494 = n3493 ^ n3431;
  assign n3495 = n3432 & ~n3494;
  assign n3496 = n3495 ^ n2583;
  assign n3497 = n3496 ^ n2374;
  assign n3498 = n3219 & ~n3397;
  assign n3499 = n3498 ^ n3241;
  assign n3500 = n3499 ^ n3496;
  assign n3501 = n3497 & ~n3500;
  assign n3502 = n3501 ^ n2374;
  assign n3503 = n3502 ^ n2194;
  assign n3504 = n3244 ^ n2374;
  assign n3505 = ~n3397 & n3504;
  assign n3506 = n3505 ^ n3246;
  assign n3507 = n3506 ^ n3502;
  assign n3508 = ~n3503 & n3507;
  assign n3509 = n3508 ^ n2194;
  assign n3510 = n3509 ^ n3416;
  assign n3511 = n3417 & n3510;
  assign n3512 = n3511 ^ n2011;
  assign n3513 = n3512 ^ n1804;
  assign n3514 = n3253 ^ n2011;
  assign n3515 = ~n3397 & ~n3514;
  assign n3516 = n3515 ^ n3182;
  assign n3517 = n3516 ^ n3512;
  assign n3518 = n3513 & n3517;
  assign n3519 = n3518 ^ n1804;
  assign n3520 = n3519 ^ n1621;
  assign n3521 = n3256 ^ n1804;
  assign n3522 = ~n3397 & n3521;
  assign n3523 = n3522 ^ n3179;
  assign n3524 = n3523 ^ n3519;
  assign n3525 = n3520 & ~n3524;
  assign n3526 = n3525 ^ n1621;
  assign n3527 = n3526 ^ n1458;
  assign n3528 = n3260 & ~n3397;
  assign n3529 = n3528 ^ n3262;
  assign n3530 = n3529 ^ n3526;
  assign n3531 = n3527 & n3530;
  assign n3532 = n3531 ^ n1458;
  assign n3533 = n3532 ^ n1299;
  assign n3534 = n3266 & ~n3397;
  assign n3535 = n3534 ^ n3269;
  assign n3536 = n3535 ^ n3532;
  assign n3537 = n3533 & ~n3536;
  assign n3538 = n3537 ^ n1299;
  assign n3539 = n3538 ^ n1158;
  assign n3540 = n3273 & ~n3397;
  assign n3541 = n3540 ^ n3276;
  assign n3542 = n3541 ^ n3538;
  assign n3543 = n3539 & ~n3542;
  assign n3544 = n3543 ^ n1158;
  assign n3545 = n3544 ^ n1027;
  assign n3546 = n3280 & ~n3397;
  assign n3547 = n3546 ^ n3282;
  assign n3548 = n3547 ^ n3544;
  assign n3549 = n3545 & ~n3548;
  assign n3550 = n3549 ^ n1027;
  assign n3551 = n3550 ^ n3412;
  assign n3552 = ~n3413 & n3551;
  assign n3553 = n3552 ^ n905;
  assign n3554 = n3553 ^ n3409;
  assign n3555 = n3410 & ~n3554;
  assign n3556 = n3555 ^ n803;
  assign n3557 = n3556 ^ n707;
  assign n3558 = n3298 & ~n3397;
  assign n3559 = n3558 ^ n3300;
  assign n3560 = n3559 ^ n3556;
  assign n3561 = ~n3557 & n3560;
  assign n3562 = n3561 ^ n707;
  assign n3563 = n3562 ^ n608;
  assign n3564 = ~n3304 & ~n3397;
  assign n3565 = n3564 ^ n3306;
  assign n3566 = n3565 ^ n3562;
  assign n3567 = ~n3563 & n3566;
  assign n3568 = n3567 ^ n608;
  assign n3571 = n3570 ^ n3568;
  assign n3572 = n3570 ^ n514;
  assign n3573 = n3571 & ~n3572;
  assign n3574 = n3573 ^ n514;
  assign n3575 = n3574 ^ n3406;
  assign n3576 = n3407 & ~n3575;
  assign n3577 = n3576 ^ n436;
  assign n3578 = n3577 ^ n363;
  assign n3579 = n3327 & ~n3397;
  assign n3580 = n3579 ^ n3329;
  assign n3581 = n3580 ^ n3577;
  assign n3582 = n3578 & n3581;
  assign n3583 = n3582 ^ n363;
  assign n3584 = n3583 ^ n300;
  assign n3585 = n3333 & ~n3397;
  assign n3586 = n3585 ^ n3335;
  assign n3587 = n3586 ^ n3583;
  assign n3588 = n3584 & ~n3587;
  assign n3589 = n3588 ^ n300;
  assign n3590 = n3404 & n3589;
  assign n3591 = n3402 ^ n210;
  assign n3592 = n243 & ~n3399;
  assign n3593 = n3592 ^ n3402;
  assign n3594 = n3591 & ~n3593;
  assign n3595 = n3594 ^ n210;
  assign n3596 = ~n3590 & ~n3595;
  assign n3597 = n3596 ^ n147;
  assign n3598 = n3353 & ~n3397;
  assign n3599 = n3598 ^ n3355;
  assign n3600 = n3599 ^ n3596;
  assign n3601 = n3597 & ~n3600;
  assign n3602 = n3601 ^ n147;
  assign n3603 = n3602 ^ n132;
  assign n3604 = ~n3359 & ~n3397;
  assign n3605 = n3604 ^ n3361;
  assign n3606 = n3605 ^ n3602;
  assign n3607 = n3603 & n3606;
  assign n3608 = n3607 ^ n132;
  assign n3619 = n1292 & n3341;
  assign n3620 = n3364 & n3619;
  assign n3609 = ~n132 & ~n3364;
  assign n3610 = n3393 & ~n3609;
  assign n3611 = n3341 & ~n3610;
  assign n3612 = ~n3341 & n3385;
  assign n3613 = n3393 & n3612;
  assign n3614 = n133 & ~n3613;
  assign n3615 = ~n3611 & n3614;
  assign n3616 = ~n133 & ~n3388;
  assign n3617 = n3393 & n3616;
  assign n3618 = ~n3615 & ~n3617;
  assign n3621 = n3620 ^ n3618;
  assign n3622 = n3621 ^ n3618;
  assign n3623 = n3618 ^ n3616;
  assign n3624 = n3623 ^ n3618;
  assign n3625 = ~n3622 & ~n3624;
  assign n3626 = n3625 ^ n3618;
  assign n3627 = n3395 & ~n3626;
  assign n3628 = n3627 ^ n3618;
  assign n3629 = n3608 & n3628;
  assign n3630 = n3385 & ~n3397;
  assign n3631 = n3630 ^ n3341;
  assign n3632 = n3628 & n3631;
  assign n3633 = ~n133 & n3632;
  assign n3634 = ~n3629 & ~n3633;
  assign n3635 = n3597 & n3634;
  assign n3636 = n3635 ^ n3599;
  assign n3637 = n3584 & n3634;
  assign n3638 = n3637 ^ n3586;
  assign n3639 = n3638 ^ n243;
  assign n3640 = n3578 & n3634;
  assign n3641 = n3640 ^ n3580;
  assign n3642 = ~n300 & n3641;
  assign n3643 = n3642 ^ n3638;
  assign n3644 = n3643 ^ n3638;
  assign n3645 = ~n3563 & n3634;
  assign n3646 = n3645 ^ n3565;
  assign n3647 = n3646 ^ n514;
  assign n3648 = ~n3557 & n3634;
  assign n3649 = n3648 ^ n3559;
  assign n3650 = n3649 ^ n608;
  assign n3651 = ~x70 & ~x71;
  assign n3652 = ~n3397 & n3651;
  assign n3653 = ~x72 & n3652;
  assign n3654 = n3634 ^ x73;
  assign n3655 = x72 & n3397;
  assign n3656 = n3397 & ~n3651;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = n3657 ^ x72;
  assign n3659 = n3658 ^ n3657;
  assign n3660 = n3657 ^ n3634;
  assign n3661 = n3660 ^ n3657;
  assign n3662 = n3659 & n3661;
  assign n3663 = n3662 ^ n3657;
  assign n3664 = n3654 & n3663;
  assign n3665 = n3664 ^ n3657;
  assign n3666 = ~n3653 & ~n3665;
  assign n3667 = n3666 ^ n3177;
  assign n3668 = n3435 ^ n3397;
  assign n3669 = n3634 & ~n3668;
  assign n3670 = n3669 ^ n3397;
  assign n3671 = n3670 ^ x74;
  assign n3672 = n3671 ^ n3666;
  assign n3673 = n3667 & n3672;
  assign n3674 = n3673 ^ n3177;
  assign n3675 = n3674 ^ n2980;
  assign n3676 = n3438 ^ n3177;
  assign n3677 = ~x74 & ~n3397;
  assign n3678 = ~n3438 & n3677;
  assign n3679 = n3676 & n3678;
  assign n3680 = n3679 ^ n3676;
  assign n3681 = n3680 ^ n3677;
  assign n3682 = n3435 ^ n3177;
  assign n3683 = n3682 ^ n3680;
  assign n3684 = n3680 ^ n3634;
  assign n3685 = ~n3680 & ~n3684;
  assign n3686 = n3685 ^ n3680;
  assign n3687 = ~n3683 & ~n3686;
  assign n3688 = n3687 ^ n3685;
  assign n3689 = n3688 ^ n3680;
  assign n3690 = n3689 ^ n3634;
  assign n3691 = n3681 & ~n3690;
  assign n3692 = n3691 ^ n3677;
  assign n3693 = n3692 ^ x75;
  assign n3694 = n3693 ^ n3674;
  assign n3695 = n3675 & ~n3694;
  assign n3696 = n3695 ^ n2980;
  assign n3697 = n3696 ^ n2782;
  assign n3708 = ~n3443 & ~n3445;
  assign n3709 = n3708 ^ x76;
  assign n3698 = x74 & ~x75;
  assign n3699 = ~n3397 & n3698;
  assign n3700 = n3436 ^ n3177;
  assign n3701 = n3397 ^ x75;
  assign n3702 = n3701 ^ n3436;
  assign n3703 = ~n3700 & n3702;
  assign n3704 = n3703 ^ n3436;
  assign n3705 = ~n3699 & ~n3704;
  assign n3706 = n3705 ^ n2980;
  assign n3707 = n3634 & n3706;
  assign n3710 = n3709 ^ n3707;
  assign n3711 = n3710 ^ n3696;
  assign n3712 = n3697 & n3711;
  assign n3713 = n3712 ^ n2782;
  assign n3714 = n3713 ^ n2583;
  assign n3715 = ~n3472 & n3634;
  assign n3716 = n3715 ^ n3490;
  assign n3717 = n3716 ^ n3713;
  assign n3718 = n3714 & ~n3717;
  assign n3719 = n3718 ^ n2583;
  assign n3720 = n3719 ^ n2374;
  assign n3721 = n3493 ^ n2583;
  assign n3722 = n3634 & n3721;
  assign n3723 = n3722 ^ n3431;
  assign n3724 = n3723 ^ n3719;
  assign n3725 = n3720 & ~n3724;
  assign n3726 = n3725 ^ n2374;
  assign n3727 = n3726 ^ n2194;
  assign n3728 = n3497 & n3634;
  assign n3729 = n3728 ^ n3499;
  assign n3730 = n3729 ^ n3726;
  assign n3731 = ~n3727 & ~n3730;
  assign n3732 = n3731 ^ n2194;
  assign n3733 = n3732 ^ n2011;
  assign n3734 = ~n3503 & n3634;
  assign n3735 = n3734 ^ n3506;
  assign n3736 = n3735 ^ n3732;
  assign n3737 = ~n3733 & ~n3736;
  assign n3738 = n3737 ^ n2011;
  assign n3739 = n3738 ^ n1804;
  assign n3740 = n3509 ^ n2011;
  assign n3741 = n3634 & ~n3740;
  assign n3742 = n3741 ^ n3416;
  assign n3743 = n3742 ^ n3738;
  assign n3744 = n3739 & ~n3743;
  assign n3745 = n3744 ^ n1804;
  assign n3746 = n3745 ^ n1621;
  assign n3747 = n3513 & n3634;
  assign n3748 = n3747 ^ n3516;
  assign n3749 = n3748 ^ n3745;
  assign n3750 = n3746 & n3749;
  assign n3751 = n3750 ^ n1621;
  assign n3752 = n3751 ^ n1458;
  assign n3753 = n3520 & n3634;
  assign n3754 = n3753 ^ n3523;
  assign n3755 = n3754 ^ n3751;
  assign n3756 = n3752 & ~n3755;
  assign n3757 = n3756 ^ n1458;
  assign n3758 = n3757 ^ n1299;
  assign n3759 = n3527 & n3634;
  assign n3760 = n3759 ^ n3529;
  assign n3761 = n3760 ^ n3757;
  assign n3762 = n3758 & n3761;
  assign n3763 = n3762 ^ n1299;
  assign n3764 = n3763 ^ n1158;
  assign n3765 = n3533 & n3634;
  assign n3766 = n3765 ^ n3535;
  assign n3767 = n3766 ^ n3763;
  assign n3768 = n3764 & ~n3767;
  assign n3769 = n3768 ^ n1158;
  assign n3770 = n3769 ^ n1027;
  assign n3771 = n3539 & n3634;
  assign n3772 = n3771 ^ n3541;
  assign n3773 = n3772 ^ n3769;
  assign n3774 = n3770 & ~n3773;
  assign n3775 = n3774 ^ n1027;
  assign n3776 = n3775 ^ n905;
  assign n3777 = n3545 & n3634;
  assign n3778 = n3777 ^ n3547;
  assign n3779 = n3778 ^ n3775;
  assign n3780 = n3776 & ~n3779;
  assign n3781 = n3780 ^ n905;
  assign n3782 = n3781 ^ n803;
  assign n3783 = n3550 ^ n905;
  assign n3784 = n3634 & n3783;
  assign n3785 = n3784 ^ n3412;
  assign n3786 = n3785 ^ n3781;
  assign n3787 = n3782 & n3786;
  assign n3788 = n3787 ^ n803;
  assign n3789 = n3788 ^ n707;
  assign n3790 = n3553 ^ n803;
  assign n3791 = n3634 & n3790;
  assign n3792 = n3791 ^ n3409;
  assign n3793 = n3792 ^ n3788;
  assign n3794 = ~n3789 & ~n3793;
  assign n3795 = n3794 ^ n707;
  assign n3796 = n3795 ^ n3649;
  assign n3797 = ~n3650 & ~n3796;
  assign n3798 = n3797 ^ n608;
  assign n3799 = n3798 ^ n3646;
  assign n3800 = n3647 & ~n3799;
  assign n3801 = n3800 ^ n514;
  assign n3802 = n436 & n3801;
  assign n3803 = n3568 ^ n514;
  assign n3804 = n3634 & n3803;
  assign n3805 = n3804 ^ n3570;
  assign n3806 = n436 & ~n3805;
  assign n3807 = ~n3802 & ~n3806;
  assign n3808 = n363 & ~n3807;
  assign n3809 = n3801 & ~n3805;
  assign n3810 = n3574 ^ n436;
  assign n3811 = n3634 & n3810;
  assign n3812 = n3811 ^ n3406;
  assign n3813 = ~n363 & ~n3812;
  assign n3814 = n3809 & ~n3813;
  assign n3815 = n436 & n3812;
  assign n3816 = n3801 & n3815;
  assign n3817 = n300 & ~n3641;
  assign n3818 = n3806 ^ n363;
  assign n3819 = n3812 ^ n3806;
  assign n3820 = ~n3806 & ~n3819;
  assign n3821 = n3820 ^ n3806;
  assign n3822 = n3818 & ~n3821;
  assign n3823 = n3822 ^ n3820;
  assign n3824 = n3823 ^ n3806;
  assign n3825 = n3824 ^ n3812;
  assign n3826 = ~n3817 & ~n3825;
  assign n3827 = n3826 ^ n3817;
  assign n3828 = ~n3816 & ~n3827;
  assign n3829 = ~n3814 & n3828;
  assign n3830 = ~n3808 & n3829;
  assign n3831 = n3830 ^ n3638;
  assign n3832 = n3831 ^ n3638;
  assign n3833 = ~n3644 & ~n3832;
  assign n3834 = n3833 ^ n3638;
  assign n3835 = n3639 & ~n3834;
  assign n3836 = n3835 ^ n243;
  assign n3837 = n3836 ^ n210;
  assign n3838 = n3589 ^ n243;
  assign n3839 = n3634 & n3838;
  assign n3840 = n3839 ^ n3399;
  assign n3841 = n3840 ^ n3836;
  assign n3842 = n3837 & n3841;
  assign n3843 = n3842 ^ n210;
  assign n3844 = n3843 ^ n147;
  assign n3845 = n3589 ^ n3399;
  assign n3846 = n3838 & n3845;
  assign n3847 = n3846 ^ n243;
  assign n3848 = n3847 ^ n210;
  assign n3849 = n3634 & n3848;
  assign n3850 = n3849 ^ n3402;
  assign n3851 = n3850 ^ n3843;
  assign n3852 = ~n3844 & ~n3851;
  assign n3853 = n3852 ^ n147;
  assign n3854 = ~n3636 & ~n3853;
  assign n3855 = n132 & ~n3854;
  assign n3856 = n3603 & n3634;
  assign n3857 = n3856 ^ n3605;
  assign n3858 = ~n133 & ~n3857;
  assign n3859 = ~n3855 & ~n3858;
  assign n3860 = n3636 & n3853;
  assign n3861 = n3859 & ~n3860;
  assign n3862 = ~n3605 & n3632;
  assign n3863 = n3608 & n3631;
  assign n3864 = n3602 & ~n3605;
  assign n3865 = ~n3628 & n3864;
  assign n3866 = ~n3631 & ~n3865;
  assign n3867 = ~n132 & n3606;
  assign n3868 = ~n3866 & ~n3867;
  assign n3869 = n3868 ^ n133;
  assign n3870 = n3869 ^ n3868;
  assign n3871 = n132 & n3602;
  assign n3872 = n3605 & ~n3871;
  assign n3873 = n3632 & n3872;
  assign n3874 = n3873 ^ n3631;
  assign n3875 = ~n3608 & ~n3874;
  assign n3876 = n3875 ^ n3868;
  assign n3877 = ~n3870 & ~n3876;
  assign n3878 = n3877 ^ n3868;
  assign n3879 = ~n3863 & n3878;
  assign n3880 = n3879 ^ n133;
  assign n3881 = ~n3862 & n3880;
  assign n3882 = ~n3861 & ~n3881;
  assign n3883 = n3651 ^ n3634;
  assign n3884 = ~n3882 & n3883;
  assign n3885 = n3884 ^ n3634;
  assign n3886 = n3885 ^ x72;
  assign n3887 = n3886 ^ n3397;
  assign n3888 = ~x68 & ~x69;
  assign n3889 = n3634 & n3888;
  assign n3890 = ~x70 & n3889;
  assign n3891 = x70 & ~n3634;
  assign n3892 = ~n3634 & ~n3888;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = n3893 ^ n3882;
  assign n3895 = n3894 ^ x71;
  assign n3896 = n3895 ^ n3882;
  assign n3897 = n3896 ^ n3894;
  assign n3898 = ~x70 & ~n3882;
  assign n3899 = n3898 ^ n3894;
  assign n3900 = ~n3897 & n3899;
  assign n3901 = n3900 ^ n3895;
  assign n3902 = ~n3890 & n3901;
  assign n3903 = n3902 ^ n3886;
  assign n3904 = n3887 & ~n3903;
  assign n3905 = n3904 ^ n3397;
  assign n3906 = n3905 ^ n3177;
  assign n3908 = n3655 ^ n3653;
  assign n3909 = n3908 ^ n3655;
  assign n3910 = n3657 ^ n3655;
  assign n3911 = n3910 ^ n3655;
  assign n3912 = ~n3909 & n3911;
  assign n3913 = n3912 ^ n3655;
  assign n3914 = ~n3634 & n3913;
  assign n3915 = n3914 ^ n3655;
  assign n3907 = ~x72 & n3634;
  assign n3916 = n3915 ^ n3907;
  assign n3917 = n3651 ^ n3397;
  assign n3918 = n3917 ^ n3915;
  assign n3919 = n3915 ^ n3882;
  assign n3920 = ~n3915 & n3919;
  assign n3921 = n3920 ^ n3915;
  assign n3922 = ~n3918 & ~n3921;
  assign n3923 = n3922 ^ n3920;
  assign n3924 = n3923 ^ n3915;
  assign n3925 = n3924 ^ n3882;
  assign n3926 = n3916 & n3925;
  assign n3927 = n3926 ^ n3907;
  assign n3928 = n3927 ^ x73;
  assign n3929 = n3928 ^ n3905;
  assign n3930 = n3906 & ~n3929;
  assign n3931 = n3930 ^ n3177;
  assign n3932 = n3931 ^ n2980;
  assign n3933 = n3667 & ~n3882;
  assign n3934 = n3933 ^ n3671;
  assign n3935 = n3934 ^ n3931;
  assign n3936 = n3932 & n3935;
  assign n3937 = n3936 ^ n2980;
  assign n3938 = n3937 ^ n2782;
  assign n3939 = n3675 & ~n3882;
  assign n3940 = n3939 ^ n3693;
  assign n3941 = n3940 ^ n3937;
  assign n3942 = n3938 & ~n3941;
  assign n3943 = n3942 ^ n2782;
  assign n3944 = n3943 ^ n2583;
  assign n3945 = n3697 & ~n3882;
  assign n3946 = n3945 ^ n3710;
  assign n3947 = n3946 ^ n3943;
  assign n3948 = n3944 & n3947;
  assign n3949 = n3948 ^ n2583;
  assign n3950 = n3949 ^ n2374;
  assign n3951 = n3714 & ~n3882;
  assign n3952 = n3951 ^ n3716;
  assign n3953 = n3952 ^ n3949;
  assign n3954 = n3950 & ~n3953;
  assign n3955 = n3954 ^ n2374;
  assign n3956 = n3955 ^ n2194;
  assign n3957 = n3720 & ~n3882;
  assign n3958 = n3957 ^ n3723;
  assign n3959 = n3958 ^ n3955;
  assign n3960 = ~n3956 & ~n3959;
  assign n3961 = n3960 ^ n2194;
  assign n3962 = n3961 ^ n2011;
  assign n3963 = ~n3727 & ~n3882;
  assign n3964 = n3963 ^ n3729;
  assign n3965 = n3964 ^ n3961;
  assign n3966 = ~n3962 & n3965;
  assign n3967 = n3966 ^ n2011;
  assign n3968 = n3967 ^ n1804;
  assign n3969 = ~n3733 & ~n3882;
  assign n3970 = n3969 ^ n3735;
  assign n3971 = n3970 ^ n3967;
  assign n3972 = n3968 & n3971;
  assign n3973 = n3972 ^ n1804;
  assign n3974 = n3973 ^ n1621;
  assign n3975 = n3739 & ~n3882;
  assign n3976 = n3975 ^ n3742;
  assign n3977 = n3976 ^ n3973;
  assign n3978 = n3974 & ~n3977;
  assign n3979 = n3978 ^ n1621;
  assign n3980 = n3979 ^ n1458;
  assign n3981 = n3746 & ~n3882;
  assign n3982 = n3981 ^ n3748;
  assign n3983 = n3982 ^ n3979;
  assign n3984 = n3980 & n3983;
  assign n3985 = n3984 ^ n1458;
  assign n3986 = n3985 ^ n1299;
  assign n3987 = n3752 & ~n3882;
  assign n3988 = n3987 ^ n3754;
  assign n3989 = n3988 ^ n3985;
  assign n3990 = n3986 & ~n3989;
  assign n3991 = n3990 ^ n1299;
  assign n3992 = n3991 ^ n1158;
  assign n3993 = n3758 & ~n3882;
  assign n3994 = n3993 ^ n3760;
  assign n3995 = n3994 ^ n3991;
  assign n3996 = n3992 & n3995;
  assign n3997 = n3996 ^ n1158;
  assign n3998 = n3997 ^ n1027;
  assign n3999 = n3853 ^ n132;
  assign n4000 = ~n3882 & n3999;
  assign n4001 = n4000 ^ n3636;
  assign n4002 = ~n133 & n4001;
  assign n4003 = n3798 ^ n514;
  assign n4004 = ~n3882 & n4003;
  assign n4005 = n4004 ^ n3646;
  assign n4006 = n4005 ^ n436;
  assign n4007 = n3795 ^ n608;
  assign n4008 = ~n3882 & ~n4007;
  assign n4009 = n4008 ^ n3649;
  assign n4010 = n4009 ^ n514;
  assign n4011 = ~n3789 & ~n3882;
  assign n4012 = n4011 ^ n3792;
  assign n4013 = ~n608 & ~n4012;
  assign n4014 = n4013 ^ n4009;
  assign n4015 = ~n4010 & n4014;
  assign n4016 = n4015 ^ n4009;
  assign n4017 = n4016 ^ n4005;
  assign n4018 = n4017 ^ n4005;
  assign n4019 = n608 & n4012;
  assign n4020 = n514 & ~n4009;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = n3776 & ~n3882;
  assign n4023 = n4022 ^ n3778;
  assign n4024 = n4023 ^ n803;
  assign n4025 = n3770 & ~n3882;
  assign n4026 = n4025 ^ n3772;
  assign n4027 = n4026 ^ n905;
  assign n4028 = n3764 & ~n3882;
  assign n4029 = n4028 ^ n3766;
  assign n4030 = n4029 ^ n3997;
  assign n4031 = n3998 & ~n4030;
  assign n4032 = n4031 ^ n1027;
  assign n4033 = n4032 ^ n4026;
  assign n4034 = n4027 & ~n4033;
  assign n4035 = n4034 ^ n905;
  assign n4036 = n4035 ^ n4023;
  assign n4037 = n4024 & ~n4036;
  assign n4038 = n4037 ^ n803;
  assign n4039 = n4038 ^ n707;
  assign n4040 = n3782 & ~n3882;
  assign n4041 = n4040 ^ n3785;
  assign n4042 = n4041 ^ n4038;
  assign n4043 = ~n4039 & n4042;
  assign n4044 = n4043 ^ n707;
  assign n4045 = n4021 & n4044;
  assign n4046 = n4045 ^ n4005;
  assign n4047 = n4046 ^ n4005;
  assign n4048 = ~n4018 & ~n4047;
  assign n4049 = n4048 ^ n4005;
  assign n4050 = n4006 & ~n4049;
  assign n4051 = n4050 ^ n436;
  assign n4052 = n4051 ^ n363;
  assign n4053 = n3801 ^ n436;
  assign n4054 = ~n3882 & n4053;
  assign n4055 = n4054 ^ n3805;
  assign n4056 = n4055 ^ n4051;
  assign n4057 = n4052 & n4056;
  assign n4058 = n4057 ^ n363;
  assign n4059 = n4058 ^ n300;
  assign n4060 = n3807 & ~n3809;
  assign n4061 = n4060 ^ n363;
  assign n4062 = ~n3882 & ~n4061;
  assign n4063 = n4062 ^ n3812;
  assign n4064 = n4063 ^ n4058;
  assign n4065 = n4059 & ~n4064;
  assign n4066 = n4065 ^ n300;
  assign n4067 = n4066 ^ n243;
  assign n4068 = n3812 ^ n363;
  assign n4069 = n4060 ^ n3812;
  assign n4070 = n4068 & n4069;
  assign n4071 = n4070 ^ n363;
  assign n4072 = n4071 ^ n300;
  assign n4073 = ~n3882 & n4072;
  assign n4074 = n4073 ^ n3641;
  assign n4075 = n4074 ^ n4066;
  assign n4076 = n4067 & n4075;
  assign n4077 = n4076 ^ n243;
  assign n4078 = n4077 ^ n210;
  assign n4079 = n3641 ^ n300;
  assign n4080 = n4071 ^ n3641;
  assign n4081 = ~n4079 & n4080;
  assign n4082 = n4081 ^ n300;
  assign n4083 = n4082 ^ n243;
  assign n4084 = ~n3882 & n4083;
  assign n4085 = n4084 ^ n3638;
  assign n4086 = n4085 ^ n4077;
  assign n4087 = n4078 & ~n4086;
  assign n4088 = n4087 ^ n210;
  assign n4089 = n4088 ^ n147;
  assign n4090 = n3837 & ~n3882;
  assign n4091 = n4090 ^ n3840;
  assign n4092 = n4091 ^ n4088;
  assign n4093 = ~n4089 & n4092;
  assign n4094 = n4093 ^ n147;
  assign n4095 = n4094 ^ n132;
  assign n4096 = ~n3844 & ~n3882;
  assign n4097 = n4096 ^ n3850;
  assign n4098 = n4097 ^ n4094;
  assign n4099 = n4095 & n4098;
  assign n4100 = n4099 ^ n132;
  assign n4101 = ~n4002 & ~n4100;
  assign n4102 = n3853 ^ n3636;
  assign n4103 = ~n3857 & n4102;
  assign n4104 = ~n132 & ~n4103;
  assign n4105 = n3857 ^ n3855;
  assign n4106 = n4105 ^ n3855;
  assign n4107 = n3860 & n3881;
  assign n4108 = n4107 ^ n3855;
  assign n4109 = n4106 & ~n4108;
  assign n4110 = n4109 ^ n3855;
  assign n4111 = n133 & ~n4110;
  assign n4112 = ~n4104 & n4111;
  assign n4113 = ~n3857 & ~n3881;
  assign n4114 = n3636 & n4113;
  assign n4115 = ~n4112 & ~n4114;
  assign n4116 = n132 & n3853;
  assign n4117 = ~n3857 & n3881;
  assign n4118 = ~n3636 & ~n4117;
  assign n4119 = ~n4116 & n4118;
  assign n4120 = n3857 ^ n132;
  assign n4121 = n4120 ^ n3853;
  assign n4122 = n4121 ^ n3857;
  assign n4123 = n3857 ^ n3853;
  assign n4124 = n4123 ^ n3853;
  assign n4125 = n4102 ^ n3853;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = n4126 ^ n3853;
  assign n4128 = n4122 & n4127;
  assign n4129 = n4128 ^ n4120;
  assign n4130 = ~n4119 & ~n4129;
  assign n4131 = ~n133 & ~n4130;
  assign n4132 = n4115 & ~n4131;
  assign n4133 = ~n4101 & ~n4132;
  assign n4134 = n3998 & ~n4133;
  assign n4135 = n4134 ^ n4029;
  assign n4136 = n4135 ^ n905;
  assign n4137 = n3992 & ~n4133;
  assign n4138 = n4137 ^ n3994;
  assign n4139 = n4138 ^ n1027;
  assign n4140 = ~x66 & ~x67;
  assign n4141 = ~n3882 & n4140;
  assign n4142 = ~x68 & n4141;
  assign n4143 = n4133 ^ x69;
  assign n4144 = x68 & n3882;
  assign n4145 = n3882 & ~n4140;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = n4146 ^ x68;
  assign n4148 = n4147 ^ n4146;
  assign n4149 = n4146 ^ n4133;
  assign n4150 = n4149 ^ n4146;
  assign n4151 = n4148 & ~n4150;
  assign n4152 = n4151 ^ n4146;
  assign n4153 = ~n4143 & n4152;
  assign n4154 = n4153 ^ n4146;
  assign n4155 = ~n4142 & ~n4154;
  assign n4156 = n4155 ^ n3634;
  assign n4157 = n3888 ^ n3882;
  assign n4158 = ~n4133 & ~n4157;
  assign n4159 = n4158 ^ n3882;
  assign n4160 = n4159 ^ x70;
  assign n4161 = n4160 ^ n4155;
  assign n4162 = ~n4156 & n4161;
  assign n4163 = n4162 ^ n3634;
  assign n4164 = n4163 ^ n3397;
  assign n4165 = ~n3890 & n3893;
  assign n4166 = n4165 ^ n3891;
  assign n4167 = n3882 & n4166;
  assign n4168 = n4167 ^ n3891;
  assign n4169 = n4168 ^ n3898;
  assign n4170 = n3888 ^ n3634;
  assign n4171 = n4170 ^ n4168;
  assign n4172 = n4168 ^ n4133;
  assign n4173 = ~n4168 & n4172;
  assign n4174 = n4173 ^ n4168;
  assign n4175 = n4171 & ~n4174;
  assign n4176 = n4175 ^ n4173;
  assign n4177 = n4176 ^ n4168;
  assign n4178 = n4177 ^ n4133;
  assign n4179 = n4169 & n4178;
  assign n4180 = n4179 ^ n3898;
  assign n4181 = n4180 ^ x71;
  assign n4182 = n4181 ^ n4163;
  assign n4183 = ~n4164 & n4182;
  assign n4184 = n4183 ^ n3397;
  assign n4185 = n4184 ^ n3177;
  assign n4186 = n3902 ^ n3397;
  assign n4187 = ~n4133 & n4186;
  assign n4188 = n4187 ^ n3886;
  assign n4189 = n4188 ^ n4184;
  assign n4190 = n4185 & ~n4189;
  assign n4191 = n4190 ^ n3177;
  assign n4192 = n4191 ^ n2980;
  assign n4193 = n3906 & ~n4133;
  assign n4194 = n4193 ^ n3928;
  assign n4195 = n4194 ^ n4191;
  assign n4196 = n4192 & ~n4195;
  assign n4197 = n4196 ^ n2980;
  assign n4198 = n4197 ^ n2782;
  assign n4199 = n3932 & ~n4133;
  assign n4200 = n4199 ^ n3934;
  assign n4201 = n4200 ^ n4197;
  assign n4202 = n4198 & n4201;
  assign n4203 = n4202 ^ n2782;
  assign n4204 = n4203 ^ n2583;
  assign n4205 = n3938 & ~n4133;
  assign n4206 = n4205 ^ n3940;
  assign n4207 = n4206 ^ n4203;
  assign n4208 = n4204 & ~n4207;
  assign n4209 = n4208 ^ n2583;
  assign n4210 = n4209 ^ n2374;
  assign n4211 = n3944 & ~n4133;
  assign n4212 = n4211 ^ n3946;
  assign n4213 = n4212 ^ n4209;
  assign n4214 = n4210 & n4213;
  assign n4215 = n4214 ^ n2374;
  assign n4216 = n4215 ^ n2194;
  assign n4217 = n3950 & ~n4133;
  assign n4218 = n4217 ^ n3952;
  assign n4219 = n4218 ^ n4215;
  assign n4220 = ~n4216 & ~n4219;
  assign n4221 = n4220 ^ n2194;
  assign n4222 = n4221 ^ n2011;
  assign n4223 = ~n3956 & ~n4133;
  assign n4224 = n4223 ^ n3958;
  assign n4225 = n4224 ^ n4221;
  assign n4226 = ~n4222 & n4225;
  assign n4227 = n4226 ^ n2011;
  assign n4228 = n4227 ^ n1804;
  assign n4229 = ~n3962 & ~n4133;
  assign n4230 = n4229 ^ n3964;
  assign n4231 = n4230 ^ n4227;
  assign n4232 = n4228 & ~n4231;
  assign n4233 = n4232 ^ n1804;
  assign n4234 = n4233 ^ n1621;
  assign n4235 = n3968 & ~n4133;
  assign n4236 = n4235 ^ n3970;
  assign n4237 = n4236 ^ n4233;
  assign n4238 = n4234 & n4237;
  assign n4239 = n4238 ^ n1621;
  assign n4240 = n4239 ^ n1458;
  assign n4241 = n3974 & ~n4133;
  assign n4242 = n4241 ^ n3976;
  assign n4243 = n4242 ^ n4239;
  assign n4244 = n4240 & ~n4243;
  assign n4245 = n4244 ^ n1458;
  assign n4246 = n4245 ^ n1299;
  assign n4247 = n3980 & ~n4133;
  assign n4248 = n4247 ^ n3982;
  assign n4249 = n4248 ^ n4245;
  assign n4250 = n4246 & n4249;
  assign n4251 = n4250 ^ n1299;
  assign n4252 = n4251 ^ n1158;
  assign n4253 = n3986 & ~n4133;
  assign n4254 = n4253 ^ n3988;
  assign n4255 = n4254 ^ n4251;
  assign n4256 = n4252 & ~n4255;
  assign n4257 = n4256 ^ n1158;
  assign n4258 = n4257 ^ n4138;
  assign n4259 = ~n4139 & n4258;
  assign n4260 = n4259 ^ n1027;
  assign n4261 = n4260 ^ n4135;
  assign n4262 = n4136 & ~n4261;
  assign n4263 = n4262 ^ n905;
  assign n4264 = n4263 ^ n803;
  assign n4265 = n133 & ~n4001;
  assign n4266 = n4101 & ~n4265;
  assign n4267 = n4115 & n4265;
  assign n4268 = ~n4002 & ~n4267;
  assign n4269 = n4100 & ~n4268;
  assign n4270 = n4001 & ~n4132;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n4266 & n4271;
  assign n4273 = ~n4089 & ~n4133;
  assign n4274 = n4273 ^ n4091;
  assign n4275 = n4274 ^ n132;
  assign n4276 = n4078 & ~n4133;
  assign n4277 = n4276 ^ n4085;
  assign n4278 = n4277 ^ n147;
  assign n4279 = n4044 ^ n608;
  assign n4280 = ~n4133 & ~n4279;
  assign n4281 = n4280 ^ n4012;
  assign n4282 = n4281 ^ n514;
  assign n4283 = ~n4039 & ~n4133;
  assign n4284 = n4283 ^ n4041;
  assign n4285 = n4284 ^ n608;
  assign n4286 = n4035 ^ n803;
  assign n4287 = ~n4133 & n4286;
  assign n4288 = n4287 ^ n4023;
  assign n4289 = n707 & ~n4288;
  assign n4290 = n4289 ^ n4284;
  assign n4291 = ~n4285 & n4290;
  assign n4292 = n4291 ^ n4284;
  assign n4293 = n4292 ^ n4281;
  assign n4294 = n4293 ^ n4281;
  assign n4295 = ~n707 & n4288;
  assign n4296 = n608 & ~n4284;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = n4032 ^ n905;
  assign n4299 = ~n4133 & n4298;
  assign n4300 = n4299 ^ n4026;
  assign n4301 = n4300 ^ n4263;
  assign n4302 = n4264 & ~n4301;
  assign n4303 = n4302 ^ n803;
  assign n4304 = n4297 & ~n4303;
  assign n4305 = n4304 ^ n4281;
  assign n4306 = n4305 ^ n4281;
  assign n4307 = ~n4294 & ~n4306;
  assign n4308 = n4307 ^ n4281;
  assign n4309 = n4282 & ~n4308;
  assign n4310 = n4309 ^ n514;
  assign n4311 = n4310 ^ n436;
  assign n4312 = n4012 ^ n608;
  assign n4313 = n4044 ^ n4012;
  assign n4314 = n4312 & n4313;
  assign n4315 = n4314 ^ n608;
  assign n4316 = n4315 ^ n514;
  assign n4317 = ~n4133 & n4316;
  assign n4318 = n4317 ^ n4009;
  assign n4319 = n4318 ^ n4310;
  assign n4320 = n4311 & n4319;
  assign n4321 = n4320 ^ n436;
  assign n4322 = n4321 ^ n363;
  assign n4323 = n4315 ^ n4009;
  assign n4324 = ~n4010 & n4323;
  assign n4325 = n4324 ^ n514;
  assign n4326 = n4325 ^ n436;
  assign n4327 = ~n4133 & n4326;
  assign n4328 = n4327 ^ n4005;
  assign n4329 = n4328 ^ n4321;
  assign n4330 = n4322 & ~n4329;
  assign n4331 = n4330 ^ n363;
  assign n4332 = n4331 ^ n300;
  assign n4333 = n4052 & ~n4133;
  assign n4334 = n4333 ^ n4055;
  assign n4335 = n4334 ^ n4331;
  assign n4336 = n4332 & n4335;
  assign n4337 = n4336 ^ n300;
  assign n4338 = n4337 ^ n243;
  assign n4339 = n4059 & ~n4133;
  assign n4340 = n4339 ^ n4063;
  assign n4341 = n4340 ^ n4337;
  assign n4342 = n4338 & ~n4341;
  assign n4343 = n4342 ^ n243;
  assign n4344 = n4343 ^ n210;
  assign n4345 = n4067 & ~n4133;
  assign n4346 = n4345 ^ n4074;
  assign n4347 = n4346 ^ n4343;
  assign n4348 = n4344 & n4347;
  assign n4349 = n4348 ^ n210;
  assign n4350 = n4349 ^ n4277;
  assign n4351 = ~n4278 & ~n4350;
  assign n4352 = n4351 ^ n147;
  assign n4353 = n4352 ^ n4274;
  assign n4354 = n4275 & ~n4353;
  assign n4355 = n4354 ^ n132;
  assign n4356 = n4355 ^ n133;
  assign n4357 = n4095 & ~n4133;
  assign n4358 = n4357 ^ n4097;
  assign n4359 = n4358 ^ n4355;
  assign n4360 = ~n4356 & ~n4359;
  assign n4361 = n4360 ^ n4355;
  assign n4362 = ~n4272 & n4361;
  assign n4363 = n4264 & ~n4362;
  assign n4364 = n4363 ^ n4300;
  assign n4365 = n4364 ^ n707;
  assign n4366 = n4260 ^ n905;
  assign n4367 = ~n4362 & n4366;
  assign n4368 = n4367 ^ n4135;
  assign n4369 = n4368 ^ n803;
  assign n4370 = n4192 & ~n4362;
  assign n4371 = n4370 ^ n4194;
  assign n4372 = n4371 ^ n2782;
  assign n4373 = n4185 & ~n4362;
  assign n4374 = n4373 ^ n4188;
  assign n4375 = n4374 ^ n2980;
  assign n4376 = ~x64 & ~x65;
  assign n4377 = ~n4133 & n4376;
  assign n4378 = ~x66 & n4377;
  assign n4379 = n4362 ^ x67;
  assign n4380 = x66 & n4133;
  assign n4381 = n4133 & ~n4376;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = n4382 ^ x66;
  assign n4384 = n4383 ^ n4382;
  assign n4385 = n4382 ^ n4362;
  assign n4386 = n4385 ^ n4382;
  assign n4387 = n4384 & ~n4386;
  assign n4388 = n4387 ^ n4382;
  assign n4389 = ~n4379 & n4388;
  assign n4390 = n4389 ^ n4382;
  assign n4391 = ~n4378 & ~n4390;
  assign n4392 = n4391 ^ n3882;
  assign n4393 = n4140 ^ n4133;
  assign n4394 = ~n4362 & ~n4393;
  assign n4395 = n4394 ^ n4133;
  assign n4396 = n4395 ^ x68;
  assign n4397 = n4396 ^ n4391;
  assign n4398 = n4392 & n4397;
  assign n4399 = n4398 ^ n3882;
  assign n4400 = n4399 ^ n3634;
  assign n4402 = n4144 ^ n4142;
  assign n4403 = n4402 ^ n4144;
  assign n4404 = n4146 ^ n4144;
  assign n4405 = n4404 ^ n4144;
  assign n4406 = ~n4403 & n4405;
  assign n4407 = n4406 ^ n4144;
  assign n4408 = n4133 & n4407;
  assign n4409 = n4408 ^ n4144;
  assign n4401 = ~x68 & ~n4133;
  assign n4410 = n4409 ^ n4401;
  assign n4411 = n4140 ^ n3882;
  assign n4412 = n4411 ^ n4409;
  assign n4413 = n4409 ^ n4362;
  assign n4414 = ~n4409 & n4413;
  assign n4415 = n4414 ^ n4409;
  assign n4416 = ~n4412 & ~n4415;
  assign n4417 = n4416 ^ n4414;
  assign n4418 = n4417 ^ n4409;
  assign n4419 = n4418 ^ n4362;
  assign n4420 = n4410 & n4419;
  assign n4421 = n4420 ^ n4401;
  assign n4422 = n4421 ^ x69;
  assign n4423 = n4422 ^ n4399;
  assign n4424 = ~n4400 & ~n4423;
  assign n4425 = n4424 ^ n3634;
  assign n4426 = n4425 ^ n3397;
  assign n4427 = ~n4156 & ~n4362;
  assign n4428 = n4427 ^ n4160;
  assign n4429 = n4428 ^ n4425;
  assign n4430 = ~n4426 & ~n4429;
  assign n4431 = n4430 ^ n3397;
  assign n4432 = n4431 ^ n3177;
  assign n4433 = ~n4164 & ~n4362;
  assign n4434 = n4433 ^ n4181;
  assign n4435 = n4434 ^ n4431;
  assign n4436 = n4432 & ~n4435;
  assign n4437 = n4436 ^ n3177;
  assign n4438 = n4437 ^ n4374;
  assign n4439 = n4375 & ~n4438;
  assign n4440 = n4439 ^ n2980;
  assign n4441 = n4440 ^ n4371;
  assign n4442 = n4372 & ~n4441;
  assign n4443 = n4442 ^ n2782;
  assign n4444 = n4443 ^ n2583;
  assign n4445 = n4198 & ~n4362;
  assign n4446 = n4445 ^ n4200;
  assign n4447 = n4446 ^ n4443;
  assign n4448 = n4444 & n4447;
  assign n4449 = n4448 ^ n2583;
  assign n4450 = n4449 ^ n2374;
  assign n4451 = n4204 & ~n4362;
  assign n4452 = n4451 ^ n4206;
  assign n4453 = n4452 ^ n4449;
  assign n4454 = n4450 & ~n4453;
  assign n4455 = n4454 ^ n2374;
  assign n4456 = n4455 ^ n2194;
  assign n4457 = n4210 & ~n4362;
  assign n4458 = n4457 ^ n4212;
  assign n4459 = n4458 ^ n4455;
  assign n4460 = ~n4456 & n4459;
  assign n4461 = n4460 ^ n2194;
  assign n4462 = n4461 ^ n2011;
  assign n4463 = ~n4216 & ~n4362;
  assign n4464 = n4463 ^ n4218;
  assign n4465 = n4464 ^ n4461;
  assign n4466 = ~n4462 & n4465;
  assign n4467 = n4466 ^ n2011;
  assign n4468 = n4467 ^ n1804;
  assign n4469 = ~n4222 & ~n4362;
  assign n4470 = n4469 ^ n4224;
  assign n4471 = n4470 ^ n4467;
  assign n4472 = n4468 & ~n4471;
  assign n4473 = n4472 ^ n1804;
  assign n4474 = n4473 ^ n1621;
  assign n4475 = n4228 & ~n4362;
  assign n4476 = n4475 ^ n4230;
  assign n4477 = n4476 ^ n4473;
  assign n4478 = n4474 & ~n4477;
  assign n4479 = n4478 ^ n1621;
  assign n4480 = n4479 ^ n1458;
  assign n4481 = n4234 & ~n4362;
  assign n4482 = n4481 ^ n4236;
  assign n4483 = n4482 ^ n4479;
  assign n4484 = n4480 & n4483;
  assign n4485 = n4484 ^ n1458;
  assign n4486 = n4485 ^ n1299;
  assign n4487 = n4240 & ~n4362;
  assign n4488 = n4487 ^ n4242;
  assign n4489 = n4488 ^ n4485;
  assign n4490 = n4486 & ~n4489;
  assign n4491 = n4490 ^ n1299;
  assign n4492 = n4491 ^ n1158;
  assign n4493 = n4246 & ~n4362;
  assign n4494 = n4493 ^ n4248;
  assign n4495 = n4494 ^ n4491;
  assign n4496 = n4492 & n4495;
  assign n4497 = n4496 ^ n1158;
  assign n4498 = n4497 ^ n1027;
  assign n4499 = n4252 & ~n4362;
  assign n4500 = n4499 ^ n4254;
  assign n4501 = n4500 ^ n4497;
  assign n4502 = n4498 & ~n4501;
  assign n4503 = n4502 ^ n1027;
  assign n4504 = n4503 ^ n905;
  assign n4505 = n4257 ^ n1027;
  assign n4506 = ~n4362 & n4505;
  assign n4507 = n4506 ^ n4138;
  assign n4508 = n4507 ^ n4503;
  assign n4509 = n4504 & n4508;
  assign n4510 = n4509 ^ n905;
  assign n4511 = n4510 ^ n4368;
  assign n4512 = n4369 & ~n4511;
  assign n4513 = n4512 ^ n803;
  assign n4514 = n4513 ^ n4364;
  assign n4515 = ~n4365 & ~n4514;
  assign n4516 = n4515 ^ n707;
  assign n4517 = n4516 ^ n608;
  assign n4518 = n4303 ^ n707;
  assign n4519 = ~n4362 & ~n4518;
  assign n4520 = n4519 ^ n4288;
  assign n4521 = n4520 ^ n4516;
  assign n4522 = ~n4517 & n4521;
  assign n4523 = n4522 ^ n608;
  assign n4524 = n4523 ^ n514;
  assign n4525 = n4288 ^ n707;
  assign n4526 = n4303 ^ n4288;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = n4527 ^ n707;
  assign n4529 = n4528 ^ n608;
  assign n4530 = ~n4362 & ~n4529;
  assign n4531 = n4530 ^ n4284;
  assign n4532 = n4531 ^ n4523;
  assign n4533 = n4524 & n4532;
  assign n4534 = n4533 ^ n514;
  assign n4535 = n4534 ^ n436;
  assign n4536 = n4528 ^ n4284;
  assign n4537 = ~n4285 & ~n4536;
  assign n4538 = n4537 ^ n608;
  assign n4539 = n4538 ^ n514;
  assign n4540 = ~n4362 & n4539;
  assign n4541 = n4540 ^ n4281;
  assign n4542 = n4541 ^ n4534;
  assign n4543 = n4535 & ~n4542;
  assign n4544 = n4543 ^ n436;
  assign n4545 = n4544 ^ n363;
  assign n4546 = n4311 & ~n4362;
  assign n4547 = n4546 ^ n4318;
  assign n4548 = n4547 ^ n4544;
  assign n4549 = n4545 & n4548;
  assign n4550 = n4549 ^ n363;
  assign n4551 = n4550 ^ n300;
  assign n4552 = n4322 & ~n4362;
  assign n4553 = n4552 ^ n4328;
  assign n4554 = n4553 ^ n4550;
  assign n4555 = n4551 & ~n4554;
  assign n4556 = n4555 ^ n300;
  assign n4557 = n4556 ^ n243;
  assign n4558 = n4332 & ~n4362;
  assign n4559 = n4558 ^ n4334;
  assign n4560 = n4559 ^ n4556;
  assign n4561 = n4557 & n4560;
  assign n4562 = n4561 ^ n243;
  assign n4563 = n4562 ^ n210;
  assign n4564 = n4338 & ~n4362;
  assign n4565 = n4564 ^ n4340;
  assign n4566 = n4565 ^ n4562;
  assign n4567 = n4563 & ~n4566;
  assign n4568 = n4567 ^ n210;
  assign n4569 = n4568 ^ n147;
  assign n4570 = n4344 & ~n4362;
  assign n4571 = n4570 ^ n4346;
  assign n4572 = n4571 ^ n4568;
  assign n4573 = ~n4569 & n4572;
  assign n4574 = n4573 ^ n147;
  assign n4575 = ~n132 & ~n4574;
  assign n4576 = n4349 ^ n147;
  assign n4577 = ~n4362 & ~n4576;
  assign n4578 = n4577 ^ n4277;
  assign n4579 = n4574 & n4578;
  assign n4580 = n132 & n4579;
  assign n4581 = n4580 ^ n4578;
  assign n4582 = ~n4575 & ~n4581;
  assign n4583 = n4352 ^ n132;
  assign n4584 = ~n4362 & n4583;
  assign n4585 = n4584 ^ n4274;
  assign n4586 = ~n133 & n4585;
  assign n4587 = ~n4582 & ~n4586;
  assign n4588 = ~n4272 & n4274;
  assign n4589 = ~n4358 & ~n4588;
  assign n4590 = n4272 ^ n133;
  assign n4591 = n4590 ^ n4272;
  assign n4592 = ~n132 & ~n4274;
  assign n4593 = ~n4352 & n4592;
  assign n4594 = n4593 ^ n4272;
  assign n4595 = n4591 & ~n4594;
  assign n4596 = n4595 ^ n4272;
  assign n4597 = ~n4355 & n4596;
  assign n4598 = n4597 ^ n133;
  assign n4599 = n4589 & n4598;
  assign n4600 = ~n133 & ~n4355;
  assign n4601 = n1292 & n4274;
  assign n4602 = n4352 & n4601;
  assign n4603 = n4358 & ~n4602;
  assign n4604 = ~n4600 & n4603;
  assign n4605 = ~n4599 & ~n4604;
  assign n4606 = ~n4587 & n4605;
  assign n4607 = n4551 & ~n4606;
  assign n4608 = n4607 ^ n4553;
  assign n4609 = ~n243 & ~n4608;
  assign n4610 = n4545 & ~n4606;
  assign n4611 = n4610 ^ n4547;
  assign n4612 = ~n300 & n4611;
  assign n4613 = ~n4609 & ~n4612;
  assign n4614 = n4376 ^ n4362;
  assign n4615 = ~n4606 & ~n4614;
  assign n4616 = n4615 ^ n4362;
  assign n4617 = n4616 ^ x66;
  assign n4618 = n4617 ^ n4133;
  assign n4619 = ~x62 & ~x63;
  assign n4620 = ~n4362 & n4619;
  assign n4621 = ~x64 & n4620;
  assign n4622 = n4606 ^ x65;
  assign n4623 = n4362 & n4619;
  assign n4624 = ~x64 & n4623;
  assign n4625 = n4624 ^ n4362;
  assign n4626 = n4625 ^ n4606;
  assign n4627 = n4626 ^ n4625;
  assign n4628 = n4625 ^ x64;
  assign n4629 = n4628 ^ n4625;
  assign n4630 = ~n4627 & n4629;
  assign n4631 = n4630 ^ n4625;
  assign n4632 = ~n4622 & ~n4631;
  assign n4633 = n4632 ^ n4625;
  assign n4634 = ~n4621 & n4633;
  assign n4635 = n4634 ^ n4617;
  assign n4636 = ~n4618 & n4635;
  assign n4637 = n4636 ^ n4133;
  assign n4638 = n4637 ^ n3882;
  assign n4640 = n4380 ^ n4378;
  assign n4641 = n4640 ^ n4380;
  assign n4642 = n4382 ^ n4380;
  assign n4643 = n4642 ^ n4380;
  assign n4644 = ~n4641 & n4643;
  assign n4645 = n4644 ^ n4380;
  assign n4646 = n4362 & n4645;
  assign n4647 = n4646 ^ n4380;
  assign n4639 = ~x66 & ~n4362;
  assign n4648 = n4647 ^ n4639;
  assign n4649 = n4376 ^ n4133;
  assign n4650 = n4649 ^ n4647;
  assign n4651 = n4647 ^ n4606;
  assign n4652 = ~n4647 & n4651;
  assign n4653 = n4652 ^ n4647;
  assign n4654 = ~n4650 & ~n4653;
  assign n4655 = n4654 ^ n4652;
  assign n4656 = n4655 ^ n4647;
  assign n4657 = n4656 ^ n4606;
  assign n4658 = n4648 & n4657;
  assign n4659 = n4658 ^ n4639;
  assign n4660 = n4659 ^ x67;
  assign n4661 = n4660 ^ n4637;
  assign n4662 = n4638 & ~n4661;
  assign n4663 = n4662 ^ n3882;
  assign n4664 = n4663 ^ n3634;
  assign n4665 = n4392 & ~n4606;
  assign n4666 = n4665 ^ n4396;
  assign n4667 = n4666 ^ n4663;
  assign n4668 = ~n4664 & n4667;
  assign n4669 = n4668 ^ n3634;
  assign n4670 = n4669 ^ n3397;
  assign n4671 = ~n4400 & ~n4606;
  assign n4672 = n4671 ^ n4422;
  assign n4673 = n4672 ^ n4669;
  assign n4674 = ~n4670 & n4673;
  assign n4675 = n4674 ^ n3397;
  assign n4676 = n4675 ^ n3177;
  assign n4677 = ~n4426 & ~n4606;
  assign n4678 = n4677 ^ n4428;
  assign n4679 = n4678 ^ n4675;
  assign n4680 = n4676 & n4679;
  assign n4681 = n4680 ^ n3177;
  assign n4682 = n4681 ^ n2980;
  assign n4683 = n4432 & ~n4606;
  assign n4684 = n4683 ^ n4434;
  assign n4685 = n4684 ^ n4681;
  assign n4686 = n4682 & ~n4685;
  assign n4687 = n4686 ^ n2980;
  assign n4688 = n4687 ^ n2782;
  assign n4689 = n4437 ^ n2980;
  assign n4690 = ~n4606 & n4689;
  assign n4691 = n4690 ^ n4374;
  assign n4692 = n4691 ^ n4687;
  assign n4693 = n4688 & ~n4692;
  assign n4694 = n4693 ^ n2782;
  assign n4695 = n4694 ^ n2583;
  assign n4696 = n4440 ^ n2782;
  assign n4697 = ~n4606 & n4696;
  assign n4698 = n4697 ^ n4371;
  assign n4699 = n4698 ^ n4694;
  assign n4700 = n4695 & ~n4699;
  assign n4701 = n4700 ^ n2583;
  assign n4702 = n4701 ^ n2374;
  assign n4703 = n4444 & ~n4606;
  assign n4704 = n4703 ^ n4446;
  assign n4705 = n4704 ^ n4701;
  assign n4706 = n4702 & n4705;
  assign n4707 = n4706 ^ n2374;
  assign n4708 = n4707 ^ n2194;
  assign n4709 = n4450 & ~n4606;
  assign n4710 = n4709 ^ n4452;
  assign n4711 = n4710 ^ n4707;
  assign n4712 = ~n4708 & ~n4711;
  assign n4713 = n4712 ^ n2194;
  assign n4714 = n4713 ^ n2011;
  assign n4715 = ~n4456 & ~n4606;
  assign n4716 = n4715 ^ n4458;
  assign n4717 = n4716 ^ n4713;
  assign n4718 = ~n4714 & ~n4717;
  assign n4719 = n4718 ^ n2011;
  assign n4720 = n4719 ^ n1804;
  assign n4721 = ~n4462 & ~n4606;
  assign n4722 = n4721 ^ n4464;
  assign n4723 = n4722 ^ n4719;
  assign n4724 = n4720 & ~n4723;
  assign n4725 = n4724 ^ n1804;
  assign n4726 = n4725 ^ n1621;
  assign n4727 = n4468 & ~n4606;
  assign n4728 = n4727 ^ n4470;
  assign n4729 = n4728 ^ n4725;
  assign n4730 = n4726 & ~n4729;
  assign n4731 = n4730 ^ n1621;
  assign n4732 = n4731 ^ n1458;
  assign n4733 = n4474 & ~n4606;
  assign n4734 = n4733 ^ n4476;
  assign n4735 = n4734 ^ n4731;
  assign n4736 = n4732 & ~n4735;
  assign n4737 = n4736 ^ n1458;
  assign n4738 = n4737 ^ n1299;
  assign n4739 = n4480 & ~n4606;
  assign n4740 = n4739 ^ n4482;
  assign n4741 = n4740 ^ n4737;
  assign n4742 = n4738 & n4741;
  assign n4743 = n4742 ^ n1299;
  assign n4744 = n4743 ^ n1158;
  assign n4745 = n4486 & ~n4606;
  assign n4746 = n4745 ^ n4488;
  assign n4747 = n4746 ^ n4743;
  assign n4748 = n4744 & ~n4747;
  assign n4749 = n4748 ^ n1158;
  assign n4750 = n4749 ^ n1027;
  assign n4751 = n4492 & ~n4606;
  assign n4752 = n4751 ^ n4494;
  assign n4753 = n4752 ^ n4749;
  assign n4754 = n4750 & n4753;
  assign n4755 = n4754 ^ n1027;
  assign n4756 = n4755 ^ n905;
  assign n4757 = n4498 & ~n4606;
  assign n4758 = n4757 ^ n4500;
  assign n4759 = n4758 ^ n4755;
  assign n4760 = n4756 & ~n4759;
  assign n4761 = n4760 ^ n905;
  assign n4762 = n4761 ^ n803;
  assign n4763 = n4504 & ~n4606;
  assign n4764 = n4763 ^ n4507;
  assign n4765 = n4764 ^ n4761;
  assign n4766 = n4762 & n4765;
  assign n4767 = n4766 ^ n803;
  assign n4768 = n4767 ^ n707;
  assign n4769 = n4510 ^ n803;
  assign n4770 = ~n4606 & n4769;
  assign n4771 = n4770 ^ n4368;
  assign n4772 = n4771 ^ n4767;
  assign n4773 = ~n4768 & ~n4772;
  assign n4774 = n4773 ^ n707;
  assign n4775 = n4774 ^ n608;
  assign n4776 = n4513 ^ n707;
  assign n4777 = ~n4606 & ~n4776;
  assign n4778 = n4777 ^ n4364;
  assign n4779 = n4778 ^ n4774;
  assign n4780 = ~n4775 & n4779;
  assign n4781 = n4780 ^ n608;
  assign n4782 = n4781 ^ n514;
  assign n4783 = ~n4517 & ~n4606;
  assign n4784 = n4783 ^ n4520;
  assign n4785 = n4784 ^ n4781;
  assign n4786 = n4782 & ~n4785;
  assign n4787 = n4786 ^ n514;
  assign n4788 = n4787 ^ n436;
  assign n4789 = n4524 & ~n4606;
  assign n4790 = n4789 ^ n4531;
  assign n4791 = n4790 ^ n4787;
  assign n4792 = n4788 & n4791;
  assign n4793 = n4792 ^ n436;
  assign n4794 = n4793 ^ n363;
  assign n4795 = n4535 & ~n4606;
  assign n4796 = n4795 ^ n4541;
  assign n4797 = n4796 ^ n4793;
  assign n4798 = n4794 & ~n4797;
  assign n4799 = n4798 ^ n363;
  assign n4800 = n4613 & n4799;
  assign n4801 = n4608 ^ n243;
  assign n4802 = n300 & ~n4611;
  assign n4803 = n4802 ^ n4608;
  assign n4804 = n4801 & ~n4803;
  assign n4805 = n4804 ^ n243;
  assign n4806 = ~n4800 & ~n4805;
  assign n4807 = n4806 ^ n210;
  assign n4808 = n4557 & ~n4606;
  assign n4809 = n4808 ^ n4559;
  assign n4810 = n4809 ^ n4806;
  assign n4811 = ~n4807 & ~n4810;
  assign n4812 = n4811 ^ n210;
  assign n4813 = n4812 ^ n147;
  assign n4814 = n4563 & ~n4606;
  assign n4815 = n4814 ^ n4565;
  assign n4816 = n4815 ^ n4812;
  assign n4817 = ~n4813 & ~n4816;
  assign n4818 = n4817 ^ n147;
  assign n4819 = n4818 ^ n132;
  assign n4820 = n4574 ^ n132;
  assign n4821 = ~n4606 & n4820;
  assign n4822 = n4821 ^ n4578;
  assign n4823 = ~n133 & ~n4822;
  assign n4824 = ~n4569 & ~n4606;
  assign n4825 = n4824 ^ n4571;
  assign n4826 = n4825 ^ n4818;
  assign n4827 = n4819 & ~n4826;
  assign n4828 = n4827 ^ n132;
  assign n4829 = ~n4823 & ~n4828;
  assign n4830 = n4582 & n4585;
  assign n4831 = n4585 & ~n4605;
  assign n4832 = n4581 & ~n4831;
  assign n4833 = n4575 & ~n4585;
  assign n4834 = ~n133 & ~n4833;
  assign n4835 = ~n4832 & n4834;
  assign n4836 = ~n4830 & n4835;
  assign n4837 = ~n4578 & n4605;
  assign n4838 = n132 & ~n4837;
  assign n4839 = n4585 ^ n4578;
  assign n4840 = n4585 ^ n4574;
  assign n4841 = ~n4839 & n4840;
  assign n4842 = n4838 & n4841;
  assign n4843 = n133 & ~n4842;
  assign n4844 = n4578 ^ n4574;
  assign n4845 = ~n132 & n4585;
  assign n4846 = ~n4844 & n4845;
  assign n4847 = n4843 & ~n4846;
  assign n4848 = ~n4836 & ~n4847;
  assign n4849 = n4585 & n4837;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4829 & ~n4850;
  assign n4852 = n4819 & ~n4851;
  assign n4853 = n4852 ^ n4825;
  assign n4854 = ~n133 & n4853;
  assign n4855 = n4794 & ~n4851;
  assign n4856 = n4855 ^ n4796;
  assign n4857 = ~n300 & ~n4856;
  assign n4858 = n4799 ^ n300;
  assign n4859 = ~n4851 & n4858;
  assign n4860 = n4859 ^ n4611;
  assign n4861 = ~n243 & n4860;
  assign n4862 = ~n4857 & ~n4861;
  assign n4863 = n4720 & ~n4851;
  assign n4864 = n4863 ^ n4722;
  assign n4865 = n4864 ^ n1621;
  assign n4866 = ~n4714 & ~n4851;
  assign n4867 = n4866 ^ n4716;
  assign n4868 = n4867 ^ n1804;
  assign n4869 = ~x60 & ~x61;
  assign n4870 = ~x62 & n4869;
  assign n4871 = n4606 & ~n4870;
  assign n4872 = n4851 ^ x63;
  assign n4873 = ~n4871 & n4872;
  assign n4875 = ~n4606 & n4869;
  assign n4874 = ~x63 & ~n4851;
  assign n4876 = n4875 ^ n4874;
  assign n4877 = ~x62 & n4876;
  assign n4878 = n4877 ^ n4874;
  assign n4879 = ~n4873 & ~n4878;
  assign n4880 = n4879 ^ n4362;
  assign n4881 = n4619 ^ n4606;
  assign n4882 = ~n4851 & ~n4881;
  assign n4883 = n4882 ^ n4606;
  assign n4884 = n4883 ^ x64;
  assign n4885 = n4884 ^ n4879;
  assign n4886 = n4880 & n4885;
  assign n4887 = n4886 ^ n4362;
  assign n4888 = n4887 ^ n4133;
  assign n4890 = n4606 ^ n4362;
  assign n4891 = n4890 ^ n4606;
  assign n4892 = n4891 ^ n4890;
  assign n4893 = n4890 ^ n4619;
  assign n4894 = n4892 & n4893;
  assign n4895 = n4894 ^ n4890;
  assign n4896 = ~x64 & n4895;
  assign n4897 = n4896 ^ n4890;
  assign n4889 = ~x64 & ~n4606;
  assign n4898 = n4897 ^ n4889;
  assign n4899 = n4619 ^ n4362;
  assign n4900 = n4899 ^ n4897;
  assign n4901 = n4897 ^ n4851;
  assign n4902 = ~n4897 & n4901;
  assign n4903 = n4902 ^ n4897;
  assign n4904 = ~n4900 & ~n4903;
  assign n4905 = n4904 ^ n4902;
  assign n4906 = n4905 ^ n4897;
  assign n4907 = n4906 ^ n4851;
  assign n4908 = n4898 & n4907;
  assign n4909 = n4908 ^ n4889;
  assign n4910 = n4909 ^ x65;
  assign n4911 = n4910 ^ n4887;
  assign n4912 = n4888 & ~n4911;
  assign n4913 = n4912 ^ n4133;
  assign n4914 = n4913 ^ n3882;
  assign n4915 = n4634 ^ n4133;
  assign n4916 = ~n4851 & n4915;
  assign n4917 = n4916 ^ n4617;
  assign n4918 = n4917 ^ n4913;
  assign n4919 = n4914 & n4918;
  assign n4920 = n4919 ^ n3882;
  assign n4921 = n4920 ^ n3634;
  assign n4922 = n4638 & ~n4851;
  assign n4923 = n4922 ^ n4660;
  assign n4924 = n4923 ^ n4920;
  assign n4925 = ~n4921 & ~n4924;
  assign n4926 = n4925 ^ n3634;
  assign n4927 = n4926 ^ n3397;
  assign n4928 = ~n4664 & ~n4851;
  assign n4929 = n4928 ^ n4666;
  assign n4930 = n4929 ^ n4926;
  assign n4931 = ~n4927 & ~n4930;
  assign n4932 = n4931 ^ n3397;
  assign n4933 = n4932 ^ n3177;
  assign n4934 = ~n4670 & ~n4851;
  assign n4935 = n4934 ^ n4672;
  assign n4936 = n4935 ^ n4932;
  assign n4937 = n4933 & ~n4936;
  assign n4938 = n4937 ^ n3177;
  assign n4939 = n4938 ^ n2980;
  assign n4940 = n4676 & ~n4851;
  assign n4941 = n4940 ^ n4678;
  assign n4942 = n4941 ^ n4938;
  assign n4943 = n4939 & n4942;
  assign n4944 = n4943 ^ n2980;
  assign n4945 = n4944 ^ n2782;
  assign n4946 = n4682 & ~n4851;
  assign n4947 = n4946 ^ n4684;
  assign n4948 = n4947 ^ n4944;
  assign n4949 = n4945 & ~n4948;
  assign n4950 = n4949 ^ n2782;
  assign n4951 = n4950 ^ n2583;
  assign n4952 = n4688 & ~n4851;
  assign n4953 = n4952 ^ n4691;
  assign n4954 = n4953 ^ n4950;
  assign n4955 = n4951 & ~n4954;
  assign n4956 = n4955 ^ n2583;
  assign n4957 = n4956 ^ n2374;
  assign n4958 = n4695 & ~n4851;
  assign n4959 = n4958 ^ n4698;
  assign n4960 = n4959 ^ n4956;
  assign n4961 = n4957 & ~n4960;
  assign n4962 = n4961 ^ n2374;
  assign n4963 = n4962 ^ n2194;
  assign n4964 = n4702 & ~n4851;
  assign n4965 = n4964 ^ n4704;
  assign n4966 = n4965 ^ n4962;
  assign n4967 = ~n4963 & n4966;
  assign n4968 = n4967 ^ n2194;
  assign n4969 = n4968 ^ n2011;
  assign n4970 = ~n4708 & ~n4851;
  assign n4971 = n4970 ^ n4710;
  assign n4972 = n4971 ^ n4968;
  assign n4973 = ~n4969 & n4972;
  assign n4974 = n4973 ^ n2011;
  assign n4975 = n4974 ^ n4867;
  assign n4976 = ~n4868 & n4975;
  assign n4977 = n4976 ^ n1804;
  assign n4978 = n4977 ^ n4864;
  assign n4979 = n4865 & ~n4978;
  assign n4980 = n4979 ^ n1621;
  assign n4981 = n1458 & n4980;
  assign n4982 = n4726 & ~n4851;
  assign n4983 = n4982 ^ n4728;
  assign n4984 = n1458 & n4983;
  assign n4985 = ~n4981 & ~n4984;
  assign n4986 = n1299 & ~n4985;
  assign n4987 = n4732 & ~n4851;
  assign n4988 = n4987 ^ n4734;
  assign n4989 = n4980 & n4983;
  assign n4990 = ~n1299 & ~n4988;
  assign n4991 = n4989 & ~n4990;
  assign n4992 = n4988 & ~n4991;
  assign n4993 = ~n1299 & ~n4984;
  assign n4994 = n4993 ^ n4991;
  assign n4995 = n4992 ^ n4981;
  assign n4996 = ~n4994 & n4995;
  assign n4997 = n4996 ^ n4981;
  assign n4998 = n4992 & n4997;
  assign n4999 = n4998 ^ n4991;
  assign n5000 = ~n4986 & ~n4999;
  assign n5001 = n5000 ^ n1158;
  assign n5002 = n4738 & ~n4851;
  assign n5003 = n5002 ^ n4740;
  assign n5004 = n5003 ^ n5000;
  assign n5005 = ~n5001 & ~n5004;
  assign n5006 = n5005 ^ n1158;
  assign n5007 = n5006 ^ n1027;
  assign n5008 = n4744 & ~n4851;
  assign n5009 = n5008 ^ n4746;
  assign n5010 = n5009 ^ n5006;
  assign n5011 = n5007 & ~n5010;
  assign n5012 = n5011 ^ n1027;
  assign n5013 = n5012 ^ n905;
  assign n5014 = n4750 & ~n4851;
  assign n5015 = n5014 ^ n4752;
  assign n5016 = n5015 ^ n5012;
  assign n5017 = n5013 & n5016;
  assign n5018 = n5017 ^ n905;
  assign n5019 = n5018 ^ n803;
  assign n5020 = n4756 & ~n4851;
  assign n5021 = n5020 ^ n4758;
  assign n5022 = n5021 ^ n5018;
  assign n5023 = n5019 & ~n5022;
  assign n5024 = n5023 ^ n803;
  assign n5025 = n5024 ^ n707;
  assign n5026 = n4762 & ~n4851;
  assign n5027 = n5026 ^ n4764;
  assign n5028 = n5027 ^ n5024;
  assign n5029 = ~n5025 & n5028;
  assign n5030 = n5029 ^ n707;
  assign n5031 = n5030 ^ n608;
  assign n5032 = ~n4768 & ~n4851;
  assign n5033 = n5032 ^ n4771;
  assign n5034 = n5033 ^ n5030;
  assign n5035 = ~n5031 & n5034;
  assign n5036 = n5035 ^ n608;
  assign n5037 = n5036 ^ n514;
  assign n5038 = ~n4775 & ~n4851;
  assign n5039 = n5038 ^ n4778;
  assign n5040 = n5039 ^ n5036;
  assign n5041 = n5037 & ~n5040;
  assign n5042 = n5041 ^ n514;
  assign n5043 = n5042 ^ n436;
  assign n5044 = n4782 & ~n4851;
  assign n5045 = n5044 ^ n4784;
  assign n5046 = n5045 ^ n5042;
  assign n5047 = n5043 & ~n5046;
  assign n5048 = n5047 ^ n436;
  assign n5049 = n5048 ^ n363;
  assign n5050 = n4788 & ~n4851;
  assign n5051 = n5050 ^ n4790;
  assign n5052 = n5051 ^ n5048;
  assign n5053 = n5049 & n5052;
  assign n5054 = n5053 ^ n363;
  assign n5055 = n4862 & n5054;
  assign n5056 = n4860 ^ n243;
  assign n5057 = n300 & n4856;
  assign n5058 = n5057 ^ n4860;
  assign n5059 = ~n5056 & n5058;
  assign n5060 = n5059 ^ n243;
  assign n5061 = ~n5055 & ~n5060;
  assign n5062 = n5061 ^ n210;
  assign n5063 = n4799 ^ n4611;
  assign n5064 = n4858 & n5063;
  assign n5065 = n5064 ^ n300;
  assign n5066 = n5065 ^ n243;
  assign n5067 = ~n4851 & n5066;
  assign n5068 = n5067 ^ n4608;
  assign n5069 = n5068 ^ n5061;
  assign n5070 = ~n5062 & n5069;
  assign n5071 = n5070 ^ n210;
  assign n5072 = n5071 ^ n147;
  assign n5073 = ~n4807 & ~n4851;
  assign n5074 = n5073 ^ n4809;
  assign n5075 = n5074 ^ n5071;
  assign n5076 = ~n5072 & n5075;
  assign n5077 = n5076 ^ n147;
  assign n5078 = n5077 ^ n132;
  assign n5079 = ~n4813 & ~n4851;
  assign n5080 = n5079 ^ n4815;
  assign n5081 = n5080 ^ n5077;
  assign n5082 = n5078 & n5081;
  assign n5083 = n5082 ^ n132;
  assign n5084 = ~n4854 & ~n5083;
  assign n5085 = ~n133 & ~n4828;
  assign n5087 = n4825 & n4850;
  assign n5088 = n1292 & n5087;
  assign n5089 = n4818 & n5088;
  assign n5090 = ~n5085 & ~n5089;
  assign n5086 = n4850 & n5085;
  assign n5091 = n5090 ^ n5086;
  assign n5092 = n5091 ^ n5090;
  assign n5093 = n4825 ^ n4819;
  assign n5094 = n5093 ^ n4850;
  assign n5095 = ~n4818 & n5087;
  assign n5096 = n5095 ^ n4850;
  assign n5097 = n5096 ^ n4850;
  assign n5098 = n5097 ^ n4825;
  assign n5099 = ~n5094 & n5098;
  assign n5100 = n5099 ^ n5093;
  assign n5101 = n133 & ~n5100;
  assign n5102 = n5101 ^ n5090;
  assign n5103 = n5102 ^ n5090;
  assign n5104 = ~n5092 & ~n5103;
  assign n5105 = n5104 ^ n5090;
  assign n5106 = ~n4822 & ~n5105;
  assign n5107 = n5106 ^ n5090;
  assign n5108 = ~n5084 & ~n5107;
  assign n5109 = n4985 & ~n4989;
  assign n5110 = n5109 ^ n1299;
  assign n5111 = ~n5108 & ~n5110;
  assign n5112 = n5111 ^ n4988;
  assign n5113 = n5112 ^ n1158;
  assign n5114 = n4980 ^ n1458;
  assign n5115 = ~n5108 & n5114;
  assign n5116 = n5115 ^ n4983;
  assign n5117 = n5116 ^ n1299;
  assign n5118 = n4914 & ~n5108;
  assign n5119 = n5118 ^ n4917;
  assign n5120 = n5119 ^ n3634;
  assign n5121 = n4888 & ~n5108;
  assign n5122 = n5121 ^ n4910;
  assign n5123 = n5122 ^ n3882;
  assign n5124 = n4869 ^ n4851;
  assign n5125 = ~n5108 & ~n5124;
  assign n5126 = n5125 ^ n4851;
  assign n5127 = n5126 ^ x62;
  assign n5128 = n5127 ^ n4606;
  assign n5129 = ~x58 & ~x59;
  assign n5130 = ~n4851 & n5129;
  assign n5131 = ~x60 & n5130;
  assign n5132 = x60 & n4851;
  assign n5133 = n4851 & ~n5129;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = n5134 ^ n5108;
  assign n5136 = n5135 ^ x61;
  assign n5137 = n5136 ^ n5108;
  assign n5138 = n5137 ^ n5135;
  assign n5139 = ~x60 & ~n5108;
  assign n5140 = n5139 ^ n5135;
  assign n5141 = ~n5138 & n5140;
  assign n5142 = n5141 ^ n5136;
  assign n5143 = ~n5131 & n5142;
  assign n5144 = n5143 ^ n5127;
  assign n5145 = ~n5128 & n5144;
  assign n5146 = n5145 ^ n4606;
  assign n5147 = n5146 ^ n4362;
  assign n5148 = ~x62 & ~n4851;
  assign n5149 = n4851 & ~n4870;
  assign n5150 = n5149 ^ n4606;
  assign n5151 = ~n5148 & n5150;
  assign n5152 = n5151 ^ n5148;
  assign n5153 = n4869 ^ n4606;
  assign n5154 = n5153 ^ n5151;
  assign n5155 = n5151 ^ n5108;
  assign n5156 = ~n5151 & n5155;
  assign n5157 = n5156 ^ n5151;
  assign n5158 = ~n5154 & ~n5157;
  assign n5159 = n5158 ^ n5156;
  assign n5160 = n5159 ^ n5151;
  assign n5161 = n5160 ^ n5108;
  assign n5162 = n5152 & n5161;
  assign n5163 = n5162 ^ n5148;
  assign n5164 = n5163 ^ x63;
  assign n5165 = n5164 ^ n5146;
  assign n5166 = n5147 & ~n5165;
  assign n5167 = n5166 ^ n4362;
  assign n5168 = n5167 ^ n4133;
  assign n5169 = n4880 & ~n5108;
  assign n5170 = n5169 ^ n4884;
  assign n5171 = n5170 ^ n5167;
  assign n5172 = n5168 & n5171;
  assign n5173 = n5172 ^ n4133;
  assign n5174 = n5173 ^ n5122;
  assign n5175 = n5123 & ~n5174;
  assign n5176 = n5175 ^ n3882;
  assign n5177 = n5176 ^ n5119;
  assign n5178 = n5120 & n5177;
  assign n5179 = n5178 ^ n3634;
  assign n5180 = n5179 ^ n3397;
  assign n5181 = ~n4921 & ~n5108;
  assign n5182 = n5181 ^ n4923;
  assign n5183 = n5182 ^ n5179;
  assign n5184 = ~n5180 & n5183;
  assign n5185 = n5184 ^ n3397;
  assign n5186 = n5185 ^ n3177;
  assign n5187 = ~n4927 & ~n5108;
  assign n5188 = n5187 ^ n4929;
  assign n5189 = n5188 ^ n5185;
  assign n5190 = n5186 & n5189;
  assign n5191 = n5190 ^ n3177;
  assign n5192 = n5191 ^ n2980;
  assign n5193 = n4933 & ~n5108;
  assign n5194 = n5193 ^ n4935;
  assign n5195 = n5194 ^ n5191;
  assign n5196 = n5192 & ~n5195;
  assign n5197 = n5196 ^ n2980;
  assign n5198 = n5197 ^ n2782;
  assign n5199 = n4939 & ~n5108;
  assign n5200 = n5199 ^ n4941;
  assign n5201 = n5200 ^ n5197;
  assign n5202 = n5198 & n5201;
  assign n5203 = n5202 ^ n2782;
  assign n5204 = n5203 ^ n2583;
  assign n5205 = n4945 & ~n5108;
  assign n5206 = n5205 ^ n4947;
  assign n5207 = n5206 ^ n5203;
  assign n5208 = n5204 & ~n5207;
  assign n5209 = n5208 ^ n2583;
  assign n5210 = n5209 ^ n2374;
  assign n5211 = n4951 & ~n5108;
  assign n5212 = n5211 ^ n4953;
  assign n5213 = n5212 ^ n5209;
  assign n5214 = n5210 & ~n5213;
  assign n5215 = n5214 ^ n2374;
  assign n5216 = n5215 ^ n2194;
  assign n5217 = n4957 & ~n5108;
  assign n5218 = n5217 ^ n4959;
  assign n5219 = n5218 ^ n5215;
  assign n5220 = ~n5216 & ~n5219;
  assign n5221 = n5220 ^ n2194;
  assign n5222 = n5221 ^ n2011;
  assign n5223 = ~n4963 & ~n5108;
  assign n5224 = n5223 ^ n4965;
  assign n5225 = n5224 ^ n5221;
  assign n5226 = ~n5222 & ~n5225;
  assign n5227 = n5226 ^ n2011;
  assign n5228 = n5227 ^ n1804;
  assign n5229 = ~n4969 & ~n5108;
  assign n5230 = n5229 ^ n4971;
  assign n5231 = n5230 ^ n5227;
  assign n5232 = n5228 & ~n5231;
  assign n5233 = n5232 ^ n1804;
  assign n5234 = n5233 ^ n1621;
  assign n5235 = n4974 ^ n1804;
  assign n5236 = ~n5108 & n5235;
  assign n5237 = n5236 ^ n4867;
  assign n5238 = n5237 ^ n5233;
  assign n5239 = n5234 & n5238;
  assign n5240 = n5239 ^ n1621;
  assign n5241 = n5240 ^ n1458;
  assign n5242 = n4977 ^ n1621;
  assign n5243 = ~n5108 & n5242;
  assign n5244 = n5243 ^ n4864;
  assign n5245 = n5244 ^ n5240;
  assign n5246 = n5241 & ~n5245;
  assign n5247 = n5246 ^ n1458;
  assign n5248 = n5247 ^ n5116;
  assign n5249 = n5117 & ~n5248;
  assign n5250 = n5249 ^ n1299;
  assign n5251 = n5250 ^ n5112;
  assign n5252 = n5113 & ~n5251;
  assign n5253 = n5252 ^ n1158;
  assign n5254 = n5253 ^ n1027;
  assign n5255 = ~n5001 & ~n5108;
  assign n5256 = n5255 ^ n5003;
  assign n5257 = n5256 ^ n5253;
  assign n5258 = n5254 & n5257;
  assign n5259 = n5258 ^ n1027;
  assign n5260 = n5259 ^ n905;
  assign n5261 = n5007 & ~n5108;
  assign n5262 = n5261 ^ n5009;
  assign n5263 = n5262 ^ n5259;
  assign n5264 = n5260 & ~n5263;
  assign n5265 = n5264 ^ n905;
  assign n5266 = n5265 ^ n803;
  assign n5267 = n5013 & ~n5108;
  assign n5268 = n5267 ^ n5015;
  assign n5269 = n5268 ^ n5265;
  assign n5270 = n5266 & n5269;
  assign n5271 = n5270 ^ n803;
  assign n5272 = n5271 ^ n707;
  assign n5273 = n5019 & ~n5108;
  assign n5274 = n5273 ^ n5021;
  assign n5275 = n5274 ^ n5271;
  assign n5276 = ~n5272 & ~n5275;
  assign n5277 = n5276 ^ n707;
  assign n5278 = n5277 ^ n608;
  assign n5279 = ~n5025 & ~n5108;
  assign n5280 = n5279 ^ n5027;
  assign n5281 = n5280 ^ n5277;
  assign n5282 = ~n5278 & ~n5281;
  assign n5283 = n5282 ^ n608;
  assign n5284 = n5283 ^ n514;
  assign n5285 = ~n5031 & ~n5108;
  assign n5286 = n5285 ^ n5033;
  assign n5287 = n5286 ^ n5283;
  assign n5288 = n5284 & ~n5287;
  assign n5289 = n5288 ^ n514;
  assign n5290 = n5289 ^ n436;
  assign n5291 = n5037 & ~n5108;
  assign n5292 = n5291 ^ n5039;
  assign n5293 = n5292 ^ n5289;
  assign n5294 = n5290 & ~n5293;
  assign n5295 = n5294 ^ n436;
  assign n5296 = n5295 ^ n363;
  assign n5297 = n5043 & ~n5108;
  assign n5298 = n5297 ^ n5045;
  assign n5299 = n5298 ^ n5295;
  assign n5300 = n5296 & ~n5299;
  assign n5301 = n5300 ^ n363;
  assign n5302 = n5301 ^ n300;
  assign n5303 = n5049 & ~n5108;
  assign n5304 = n5303 ^ n5051;
  assign n5305 = n5304 ^ n5301;
  assign n5306 = n5302 & n5305;
  assign n5307 = n5306 ^ n300;
  assign n5308 = n5307 ^ n243;
  assign n5309 = n5054 ^ n300;
  assign n5310 = ~n5108 & n5309;
  assign n5311 = n5310 ^ n4856;
  assign n5312 = n5311 ^ n5307;
  assign n5313 = n5308 & ~n5312;
  assign n5314 = n5313 ^ n243;
  assign n5315 = n5314 ^ n210;
  assign n5316 = n5054 ^ n4856;
  assign n5317 = n5309 & ~n5316;
  assign n5318 = n5317 ^ n300;
  assign n5319 = n5318 ^ n243;
  assign n5320 = ~n5108 & n5319;
  assign n5321 = n5320 ^ n4860;
  assign n5322 = n5321 ^ n5314;
  assign n5323 = n5315 & n5322;
  assign n5324 = n5323 ^ n210;
  assign n5325 = n5324 ^ n147;
  assign n5326 = ~n5062 & ~n5108;
  assign n5327 = n5326 ^ n5068;
  assign n5328 = n5327 ^ n5324;
  assign n5329 = ~n5325 & ~n5328;
  assign n5330 = n5329 ^ n147;
  assign n5331 = n5330 ^ n132;
  assign n5332 = ~n132 & ~n5077;
  assign n5333 = n5332 ^ n5080;
  assign n5334 = n132 & n5077;
  assign n5335 = ~n5108 & ~n5334;
  assign n5336 = ~n5332 & ~n5335;
  assign n5337 = n5333 & n5336;
  assign n5338 = n5337 ^ n5333;
  assign n5339 = n4853 & n5338;
  assign n5340 = n5108 & ~n5332;
  assign n5341 = ~n4853 & n5334;
  assign n5342 = ~n5340 & ~n5341;
  assign n5343 = ~n5080 & ~n5342;
  assign n5344 = ~n5339 & ~n5343;
  assign n5345 = ~n5072 & ~n5108;
  assign n5346 = n5345 ^ n5074;
  assign n5347 = n5346 ^ n5330;
  assign n5348 = n5331 & ~n5347;
  assign n5349 = n5348 ^ n132;
  assign n5350 = ~n5344 & n5349;
  assign n5351 = n133 & ~n5350;
  assign n5352 = ~n5332 & n5335;
  assign n5353 = n5352 ^ n5080;
  assign n5354 = ~n5349 & n5353;
  assign n5355 = n5083 ^ n4853;
  assign n5356 = n4853 ^ n133;
  assign n5357 = n5107 ^ n133;
  assign n5358 = n5357 ^ n133;
  assign n5359 = n5356 & ~n5358;
  assign n5360 = n5359 ^ n133;
  assign n5361 = n5355 & ~n5360;
  assign n5362 = ~n5354 & ~n5361;
  assign n5363 = ~n5351 & n5362;
  assign n5364 = n5331 & ~n5363;
  assign n5365 = n5364 ^ n5346;
  assign n5366 = ~n133 & n5365;
  assign n5367 = n5302 & ~n5363;
  assign n5368 = n5367 ^ n5304;
  assign n5369 = ~n243 & n5368;
  assign n5370 = n5308 & ~n5363;
  assign n5371 = n5370 ^ n5311;
  assign n5372 = ~n210 & ~n5371;
  assign n5373 = ~n5369 & ~n5372;
  assign n5374 = n5290 & ~n5363;
  assign n5375 = n5374 ^ n5292;
  assign n5376 = n5375 ^ n363;
  assign n5377 = n5284 & ~n5363;
  assign n5378 = n5377 ^ n5286;
  assign n5379 = n5378 ^ n436;
  assign n5380 = n5241 & ~n5363;
  assign n5381 = n5380 ^ n5244;
  assign n5382 = n5381 ^ n1299;
  assign n5383 = n5234 & ~n5363;
  assign n5384 = n5383 ^ n5237;
  assign n5385 = n5384 ^ n1458;
  assign n5386 = n5198 & ~n5363;
  assign n5387 = n5386 ^ n5200;
  assign n5388 = n5387 ^ n2583;
  assign n5389 = n5192 & ~n5363;
  assign n5390 = n5389 ^ n5194;
  assign n5391 = n5390 ^ n2782;
  assign n5392 = n5129 ^ n5108;
  assign n5393 = ~n5363 & ~n5392;
  assign n5394 = n5393 ^ n5108;
  assign n5395 = n5394 ^ x60;
  assign n5396 = n5395 ^ n4851;
  assign n5397 = ~x56 & ~x57;
  assign n5398 = ~n5108 & n5397;
  assign n5399 = ~x58 & n5398;
  assign n5400 = n5363 ^ x59;
  assign n5401 = n5108 & n5397;
  assign n5402 = ~x58 & n5401;
  assign n5403 = n5402 ^ n5108;
  assign n5404 = n5403 ^ n5363;
  assign n5405 = n5404 ^ n5403;
  assign n5406 = n5403 ^ x58;
  assign n5407 = n5406 ^ n5403;
  assign n5408 = ~n5405 & n5407;
  assign n5409 = n5408 ^ n5403;
  assign n5410 = ~n5400 & ~n5409;
  assign n5411 = n5410 ^ n5403;
  assign n5412 = ~n5399 & n5411;
  assign n5413 = n5412 ^ n5395;
  assign n5414 = ~n5396 & n5413;
  assign n5415 = n5414 ^ n4851;
  assign n5416 = n5415 ^ n4606;
  assign n5417 = ~n5131 & n5134;
  assign n5418 = n5417 ^ n5132;
  assign n5419 = n5108 & n5418;
  assign n5420 = n5419 ^ n5132;
  assign n5421 = n5420 ^ n5139;
  assign n5422 = n5129 ^ n4851;
  assign n5423 = n5422 ^ n5420;
  assign n5424 = n5420 ^ n5363;
  assign n5425 = ~n5420 & n5424;
  assign n5426 = n5425 ^ n5420;
  assign n5427 = ~n5423 & ~n5426;
  assign n5428 = n5427 ^ n5425;
  assign n5429 = n5428 ^ n5420;
  assign n5430 = n5429 ^ n5363;
  assign n5431 = n5421 & n5430;
  assign n5432 = n5431 ^ n5139;
  assign n5433 = n5432 ^ x61;
  assign n5434 = n5433 ^ n5415;
  assign n5435 = n5416 & ~n5434;
  assign n5436 = n5435 ^ n4606;
  assign n5437 = n5436 ^ n4362;
  assign n5438 = n5143 ^ n4606;
  assign n5439 = ~n5363 & n5438;
  assign n5440 = n5439 ^ n5127;
  assign n5441 = n5440 ^ n5436;
  assign n5442 = n5437 & n5441;
  assign n5443 = n5442 ^ n4362;
  assign n5444 = n5443 ^ n4133;
  assign n5445 = n5147 & ~n5363;
  assign n5446 = n5445 ^ n5164;
  assign n5447 = n5446 ^ n5443;
  assign n5448 = n5444 & ~n5447;
  assign n5449 = n5448 ^ n4133;
  assign n5450 = n5449 ^ n3882;
  assign n5451 = n5168 & ~n5363;
  assign n5452 = n5451 ^ n5170;
  assign n5453 = n5452 ^ n5449;
  assign n5454 = n5450 & n5453;
  assign n5455 = n5454 ^ n3882;
  assign n5456 = n5455 ^ n3634;
  assign n5457 = n5173 ^ n3882;
  assign n5458 = ~n5363 & n5457;
  assign n5459 = n5458 ^ n5122;
  assign n5460 = n5459 ^ n5455;
  assign n5461 = ~n5456 & ~n5460;
  assign n5462 = n5461 ^ n3634;
  assign n5463 = n5462 ^ n3397;
  assign n5464 = n5176 ^ n3634;
  assign n5465 = ~n5363 & ~n5464;
  assign n5466 = n5465 ^ n5119;
  assign n5467 = n5466 ^ n5462;
  assign n5468 = ~n5463 & ~n5467;
  assign n5469 = n5468 ^ n3397;
  assign n5470 = n5469 ^ n3177;
  assign n5471 = ~n5180 & ~n5363;
  assign n5472 = n5471 ^ n5182;
  assign n5473 = n5472 ^ n5469;
  assign n5474 = n5470 & ~n5473;
  assign n5475 = n5474 ^ n3177;
  assign n5476 = n5475 ^ n2980;
  assign n5477 = n5186 & ~n5363;
  assign n5478 = n5477 ^ n5188;
  assign n5479 = n5478 ^ n5475;
  assign n5480 = n5476 & n5479;
  assign n5481 = n5480 ^ n2980;
  assign n5482 = n5481 ^ n5390;
  assign n5483 = n5391 & ~n5482;
  assign n5484 = n5483 ^ n2782;
  assign n5485 = n5484 ^ n5387;
  assign n5486 = ~n5388 & n5485;
  assign n5487 = n5486 ^ n2583;
  assign n5488 = n5487 ^ n2374;
  assign n5489 = n5204 & ~n5363;
  assign n5490 = n5489 ^ n5206;
  assign n5491 = n5490 ^ n5487;
  assign n5492 = n5488 & ~n5491;
  assign n5493 = n5492 ^ n2374;
  assign n5494 = n5493 ^ n2194;
  assign n5495 = n5210 & ~n5363;
  assign n5496 = n5495 ^ n5212;
  assign n5497 = n5496 ^ n5493;
  assign n5498 = ~n5494 & ~n5497;
  assign n5499 = n5498 ^ n2194;
  assign n5500 = n5499 ^ n2011;
  assign n5501 = ~n5216 & ~n5363;
  assign n5502 = n5501 ^ n5218;
  assign n5503 = n5502 ^ n5499;
  assign n5504 = ~n5500 & n5503;
  assign n5505 = n5504 ^ n2011;
  assign n5506 = n5505 ^ n1804;
  assign n5507 = ~n5222 & ~n5363;
  assign n5508 = n5507 ^ n5224;
  assign n5509 = n5508 ^ n5505;
  assign n5510 = n5506 & n5509;
  assign n5511 = n5510 ^ n1804;
  assign n5512 = n5511 ^ n1621;
  assign n5513 = n5228 & ~n5363;
  assign n5514 = n5513 ^ n5230;
  assign n5515 = n5514 ^ n5511;
  assign n5516 = n5512 & ~n5515;
  assign n5517 = n5516 ^ n1621;
  assign n5518 = n5517 ^ n5384;
  assign n5519 = ~n5385 & n5518;
  assign n5520 = n5519 ^ n1458;
  assign n5521 = n5520 ^ n5381;
  assign n5522 = n5382 & ~n5521;
  assign n5523 = n5522 ^ n1299;
  assign n5524 = n5523 ^ n1158;
  assign n5525 = n5247 ^ n1299;
  assign n5526 = ~n5363 & n5525;
  assign n5527 = n5526 ^ n5116;
  assign n5528 = n5527 ^ n5523;
  assign n5529 = n5524 & ~n5528;
  assign n5530 = n5529 ^ n1158;
  assign n5531 = n5530 ^ n1027;
  assign n5532 = n5250 ^ n1158;
  assign n5533 = ~n5363 & n5532;
  assign n5534 = n5533 ^ n5112;
  assign n5535 = n5534 ^ n5530;
  assign n5536 = n5531 & ~n5535;
  assign n5537 = n5536 ^ n1027;
  assign n5538 = n5537 ^ n905;
  assign n5539 = n5254 & ~n5363;
  assign n5540 = n5539 ^ n5256;
  assign n5541 = n5540 ^ n5537;
  assign n5542 = n5538 & n5541;
  assign n5543 = n5542 ^ n905;
  assign n5544 = n5543 ^ n803;
  assign n5545 = n5260 & ~n5363;
  assign n5546 = n5545 ^ n5262;
  assign n5547 = n5546 ^ n5543;
  assign n5548 = n5544 & ~n5547;
  assign n5549 = n5548 ^ n803;
  assign n5550 = n5549 ^ n707;
  assign n5551 = n5266 & ~n5363;
  assign n5552 = n5551 ^ n5268;
  assign n5553 = n5552 ^ n5549;
  assign n5554 = ~n5550 & n5553;
  assign n5555 = n5554 ^ n707;
  assign n5556 = n5555 ^ n608;
  assign n5557 = ~n5272 & ~n5363;
  assign n5558 = n5557 ^ n5274;
  assign n5559 = n5558 ^ n5555;
  assign n5560 = ~n5556 & n5559;
  assign n5561 = n5560 ^ n608;
  assign n5562 = n5561 ^ n514;
  assign n5563 = ~n5278 & ~n5363;
  assign n5564 = n5563 ^ n5280;
  assign n5565 = n5564 ^ n5561;
  assign n5566 = n5562 & n5565;
  assign n5567 = n5566 ^ n514;
  assign n5568 = n5567 ^ n5378;
  assign n5569 = n5379 & ~n5568;
  assign n5570 = n5569 ^ n436;
  assign n5571 = n5570 ^ n5375;
  assign n5572 = n5376 & ~n5571;
  assign n5573 = n5572 ^ n363;
  assign n5574 = n5573 ^ n300;
  assign n5575 = n5296 & ~n5363;
  assign n5576 = n5575 ^ n5298;
  assign n5577 = n5576 ^ n5573;
  assign n5578 = n5574 & ~n5577;
  assign n5579 = n5578 ^ n300;
  assign n5580 = n5373 & n5579;
  assign n5581 = n5371 ^ n210;
  assign n5582 = n243 & ~n5368;
  assign n5583 = n5582 ^ n5371;
  assign n5584 = n5581 & ~n5583;
  assign n5585 = n5584 ^ n210;
  assign n5586 = ~n5580 & ~n5585;
  assign n5587 = n5586 ^ n147;
  assign n5588 = n5315 & ~n5363;
  assign n5589 = n5588 ^ n5321;
  assign n5590 = n5589 ^ n5586;
  assign n5591 = n5587 & ~n5590;
  assign n5592 = n5591 ^ n147;
  assign n5593 = n5592 ^ n132;
  assign n5594 = ~n5325 & ~n5363;
  assign n5595 = n5594 ^ n5327;
  assign n5596 = n5595 ^ n5592;
  assign n5597 = n5593 & n5596;
  assign n5598 = n5597 ^ n132;
  assign n5599 = ~n5366 & ~n5598;
  assign n5601 = ~n5330 & ~n5346;
  assign n5609 = x127 & n5601;
  assign n5610 = n5330 & n5346;
  assign n5611 = n5610 ^ n1292;
  assign n5612 = n5611 ^ n1292;
  assign n5613 = n130 ^ x127;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = n5614 ^ n1292;
  assign n5616 = ~n5609 & ~n5615;
  assign n5600 = n5346 & n5363;
  assign n5602 = ~n132 & n5601;
  assign n5603 = n133 & ~n5602;
  assign n5604 = ~n5349 & n5603;
  assign n5605 = ~n5600 & ~n5604;
  assign n5606 = ~n5349 & ~n5362;
  assign n5607 = ~n133 & ~n5606;
  assign n5608 = n5605 & ~n5607;
  assign n5617 = n5616 ^ n5608;
  assign n5618 = n5617 ^ n5608;
  assign n5619 = n5608 ^ n5363;
  assign n5620 = n5619 ^ n5608;
  assign n5621 = ~n5618 & ~n5620;
  assign n5622 = n5621 ^ n5608;
  assign n5623 = n5353 & ~n5622;
  assign n5624 = n5623 ^ n5608;
  assign n5625 = ~n5599 & ~n5624;
  assign n5626 = n5570 ^ n363;
  assign n5627 = ~n5625 & n5626;
  assign n5628 = n5627 ^ n5375;
  assign n5629 = n5628 ^ n300;
  assign n5630 = n5567 ^ n436;
  assign n5631 = ~n5625 & n5630;
  assign n5632 = n5631 ^ n5378;
  assign n5633 = n5632 ^ n363;
  assign n5634 = n5538 & ~n5625;
  assign n5635 = n5634 ^ n5540;
  assign n5636 = n5635 ^ n803;
  assign n5637 = n5531 & ~n5625;
  assign n5638 = n5637 ^ n5534;
  assign n5639 = n5638 ^ n905;
  assign n5640 = n5484 ^ n2583;
  assign n5641 = ~n5625 & n5640;
  assign n5642 = n5641 ^ n5387;
  assign n5643 = n5642 ^ n2374;
  assign n5644 = n5481 ^ n2782;
  assign n5645 = ~n5625 & n5644;
  assign n5646 = n5645 ^ n5390;
  assign n5647 = n5646 ^ n2583;
  assign n5648 = ~x54 & ~x55;
  assign n5649 = ~n5363 & n5648;
  assign n5650 = ~x56 & n5649;
  assign n5651 = n5625 ^ x57;
  assign n5652 = x56 & n5363;
  assign n5653 = n5363 & ~n5648;
  assign n5654 = ~n5652 & ~n5653;
  assign n5655 = n5654 ^ x56;
  assign n5656 = n5655 ^ n5654;
  assign n5657 = n5654 ^ n5625;
  assign n5658 = n5657 ^ n5654;
  assign n5659 = n5656 & ~n5658;
  assign n5660 = n5659 ^ n5654;
  assign n5661 = ~n5651 & n5660;
  assign n5662 = n5661 ^ n5654;
  assign n5663 = ~n5650 & ~n5662;
  assign n5664 = n5663 ^ n5108;
  assign n5665 = n5397 ^ n5363;
  assign n5666 = ~n5625 & ~n5665;
  assign n5667 = n5666 ^ n5363;
  assign n5668 = n5667 ^ x58;
  assign n5669 = n5668 ^ n5663;
  assign n5670 = n5664 & n5669;
  assign n5671 = n5670 ^ n5108;
  assign n5672 = n5671 ^ n4851;
  assign n5674 = n5363 ^ n5108;
  assign n5675 = n5674 ^ n5363;
  assign n5676 = n5675 ^ n5674;
  assign n5677 = n5674 ^ n5397;
  assign n5678 = n5676 & n5677;
  assign n5679 = n5678 ^ n5674;
  assign n5680 = ~x58 & n5679;
  assign n5681 = n5680 ^ n5674;
  assign n5673 = ~x58 & ~n5363;
  assign n5682 = n5681 ^ n5673;
  assign n5683 = n5397 ^ n5108;
  assign n5684 = n5683 ^ n5681;
  assign n5685 = n5681 ^ n5625;
  assign n5686 = ~n5681 & n5685;
  assign n5687 = n5686 ^ n5681;
  assign n5688 = ~n5684 & ~n5687;
  assign n5689 = n5688 ^ n5686;
  assign n5690 = n5689 ^ n5681;
  assign n5691 = n5690 ^ n5625;
  assign n5692 = n5682 & n5691;
  assign n5693 = n5692 ^ n5673;
  assign n5694 = n5693 ^ x59;
  assign n5695 = n5694 ^ n5671;
  assign n5696 = n5672 & ~n5695;
  assign n5697 = n5696 ^ n4851;
  assign n5698 = n5697 ^ n4606;
  assign n5699 = n5412 ^ n4851;
  assign n5700 = ~n5625 & n5699;
  assign n5701 = n5700 ^ n5395;
  assign n5702 = n5701 ^ n5697;
  assign n5703 = n5698 & n5702;
  assign n5704 = n5703 ^ n4606;
  assign n5705 = n5704 ^ n4362;
  assign n5706 = n5416 & ~n5625;
  assign n5707 = n5706 ^ n5433;
  assign n5708 = n5707 ^ n5704;
  assign n5709 = n5705 & ~n5708;
  assign n5710 = n5709 ^ n4362;
  assign n5711 = n5710 ^ n4133;
  assign n5712 = n5437 & ~n5625;
  assign n5713 = n5712 ^ n5440;
  assign n5714 = n5713 ^ n5710;
  assign n5715 = n5711 & n5714;
  assign n5716 = n5715 ^ n4133;
  assign n5717 = n5716 ^ n3882;
  assign n5718 = n5444 & ~n5625;
  assign n5719 = n5718 ^ n5446;
  assign n5720 = n5719 ^ n5716;
  assign n5721 = n5717 & ~n5720;
  assign n5722 = n5721 ^ n3882;
  assign n5723 = n5722 ^ n3634;
  assign n5724 = n5450 & ~n5625;
  assign n5725 = n5724 ^ n5452;
  assign n5726 = n5725 ^ n5722;
  assign n5727 = ~n5723 & n5726;
  assign n5728 = n5727 ^ n3634;
  assign n5729 = n5728 ^ n3397;
  assign n5730 = ~n5456 & ~n5625;
  assign n5731 = n5730 ^ n5459;
  assign n5732 = n5731 ^ n5728;
  assign n5733 = ~n5729 & n5732;
  assign n5734 = n5733 ^ n3397;
  assign n5735 = n5734 ^ n3177;
  assign n5736 = ~n5463 & ~n5625;
  assign n5737 = n5736 ^ n5466;
  assign n5738 = n5737 ^ n5734;
  assign n5739 = n5735 & n5738;
  assign n5740 = n5739 ^ n3177;
  assign n5741 = n5740 ^ n2980;
  assign n5742 = n5470 & ~n5625;
  assign n5743 = n5742 ^ n5472;
  assign n5744 = n5743 ^ n5740;
  assign n5745 = n5741 & ~n5744;
  assign n5746 = n5745 ^ n2980;
  assign n5747 = n5746 ^ n2782;
  assign n5748 = n5476 & ~n5625;
  assign n5749 = n5748 ^ n5478;
  assign n5750 = n5749 ^ n5746;
  assign n5751 = n5747 & n5750;
  assign n5752 = n5751 ^ n2782;
  assign n5753 = n5752 ^ n5646;
  assign n5754 = n5647 & ~n5753;
  assign n5755 = n5754 ^ n2583;
  assign n5756 = n5755 ^ n5642;
  assign n5757 = ~n5643 & n5756;
  assign n5758 = n5757 ^ n2374;
  assign n5759 = n5758 ^ n2194;
  assign n5760 = n5488 & ~n5625;
  assign n5761 = n5760 ^ n5490;
  assign n5762 = n5761 ^ n5758;
  assign n5763 = ~n5759 & ~n5762;
  assign n5764 = n5763 ^ n2194;
  assign n5765 = n5764 ^ n2011;
  assign n5766 = ~n5494 & ~n5625;
  assign n5767 = n5766 ^ n5496;
  assign n5768 = n5767 ^ n5764;
  assign n5769 = ~n5765 & n5768;
  assign n5770 = n5769 ^ n2011;
  assign n5771 = n5770 ^ n1804;
  assign n5772 = ~n5500 & ~n5625;
  assign n5773 = n5772 ^ n5502;
  assign n5774 = n5773 ^ n5770;
  assign n5775 = n5771 & ~n5774;
  assign n5776 = n5775 ^ n1804;
  assign n5777 = n5776 ^ n1621;
  assign n5778 = n5506 & ~n5625;
  assign n5779 = n5778 ^ n5508;
  assign n5780 = n5779 ^ n5776;
  assign n5781 = n5777 & n5780;
  assign n5782 = n5781 ^ n1621;
  assign n5783 = n5782 ^ n1458;
  assign n5784 = n5512 & ~n5625;
  assign n5785 = n5784 ^ n5514;
  assign n5786 = n5785 ^ n5782;
  assign n5787 = n5783 & ~n5786;
  assign n5788 = n5787 ^ n1458;
  assign n5789 = n5788 ^ n1299;
  assign n5790 = n5517 ^ n1458;
  assign n5791 = ~n5625 & n5790;
  assign n5792 = n5791 ^ n5384;
  assign n5793 = n5792 ^ n5788;
  assign n5794 = n5789 & n5793;
  assign n5795 = n5794 ^ n1299;
  assign n5796 = n5795 ^ n1158;
  assign n5797 = n5520 ^ n1299;
  assign n5798 = ~n5625 & n5797;
  assign n5799 = n5798 ^ n5381;
  assign n5800 = n5799 ^ n5795;
  assign n5801 = n5796 & ~n5800;
  assign n5802 = n5801 ^ n1158;
  assign n5803 = n5802 ^ n1027;
  assign n5804 = n5524 & ~n5625;
  assign n5805 = n5804 ^ n5527;
  assign n5806 = n5805 ^ n5802;
  assign n5807 = n5803 & ~n5806;
  assign n5808 = n5807 ^ n1027;
  assign n5809 = n5808 ^ n5638;
  assign n5810 = n5639 & ~n5809;
  assign n5811 = n5810 ^ n905;
  assign n5812 = n5811 ^ n5635;
  assign n5813 = ~n5636 & n5812;
  assign n5814 = n5813 ^ n803;
  assign n5815 = n5814 ^ n707;
  assign n5816 = n5544 & ~n5625;
  assign n5817 = n5816 ^ n5546;
  assign n5818 = n5817 ^ n5814;
  assign n5819 = ~n5815 & ~n5818;
  assign n5820 = n5819 ^ n707;
  assign n5821 = n5820 ^ n608;
  assign n5822 = ~n5550 & ~n5625;
  assign n5823 = n5822 ^ n5552;
  assign n5824 = n5823 ^ n5820;
  assign n5825 = ~n5821 & ~n5824;
  assign n5826 = n5825 ^ n608;
  assign n5827 = n5826 ^ n514;
  assign n5828 = ~n5556 & ~n5625;
  assign n5829 = n5828 ^ n5558;
  assign n5830 = n5829 ^ n5826;
  assign n5831 = n5827 & ~n5830;
  assign n5832 = n5831 ^ n514;
  assign n5833 = n5832 ^ n436;
  assign n5834 = n5562 & ~n5625;
  assign n5835 = n5834 ^ n5564;
  assign n5836 = n5835 ^ n5832;
  assign n5837 = n5833 & n5836;
  assign n5838 = n5837 ^ n436;
  assign n5839 = n5838 ^ n5632;
  assign n5840 = n5633 & ~n5839;
  assign n5841 = n5840 ^ n363;
  assign n5842 = n5841 ^ n5628;
  assign n5843 = n5629 & ~n5842;
  assign n5844 = n5843 ^ n300;
  assign n5845 = n5844 ^ n243;
  assign n5846 = n5574 & ~n5625;
  assign n5847 = n5846 ^ n5576;
  assign n5848 = n5847 ^ n5844;
  assign n5849 = n5845 & ~n5848;
  assign n5850 = n5849 ^ n243;
  assign n5851 = n5850 ^ n210;
  assign n5852 = n5579 ^ n243;
  assign n5853 = ~n5625 & n5852;
  assign n5854 = n5853 ^ n5368;
  assign n5855 = n5854 ^ n5850;
  assign n5856 = n5851 & n5855;
  assign n5857 = n5856 ^ n210;
  assign n5858 = n5857 ^ n147;
  assign n5859 = n5593 & ~n5625;
  assign n5860 = n5859 ^ n5595;
  assign n5861 = ~n133 & ~n5860;
  assign n5862 = n5579 ^ n5368;
  assign n5863 = n5852 & n5862;
  assign n5864 = n5863 ^ n243;
  assign n5865 = n5864 ^ n210;
  assign n5866 = ~n5625 & n5865;
  assign n5867 = n5866 ^ n5371;
  assign n5868 = n5867 ^ n5857;
  assign n5869 = ~n5858 & ~n5868;
  assign n5870 = n5869 ^ n147;
  assign n5871 = n5870 ^ n132;
  assign n5872 = n5587 & ~n5625;
  assign n5873 = n5872 ^ n5589;
  assign n5874 = n5873 ^ n5870;
  assign n5875 = n5871 & ~n5874;
  assign n5876 = n5875 ^ n132;
  assign n5877 = ~n5861 & ~n5876;
  assign n5878 = n133 & n5365;
  assign n5879 = n5595 ^ n5593;
  assign n5880 = n5879 ^ n5624;
  assign n5881 = ~n5595 & n5624;
  assign n5882 = ~n5592 & n5881;
  assign n5883 = n5882 ^ n5624;
  assign n5884 = n5883 ^ n5624;
  assign n5885 = n5884 ^ n5595;
  assign n5886 = n5880 & ~n5885;
  assign n5887 = n5886 ^ n5879;
  assign n5888 = n5878 & n5887;
  assign n5892 = n5366 & n5624;
  assign n5889 = n1292 & n5881;
  assign n5890 = n5592 & n5889;
  assign n5891 = ~n5365 & ~n5890;
  assign n5893 = n5892 ^ n5891;
  assign n5894 = n5892 ^ n133;
  assign n5895 = n5892 ^ n5598;
  assign n5896 = ~n5892 & n5895;
  assign n5897 = n5896 ^ n5892;
  assign n5898 = ~n5894 & ~n5897;
  assign n5899 = n5898 ^ n5896;
  assign n5900 = n5899 ^ n5892;
  assign n5901 = n5900 ^ n5598;
  assign n5902 = n5893 & n5901;
  assign n5903 = n5902 ^ n5891;
  assign n5904 = ~n5888 & ~n5903;
  assign n5905 = ~n5877 & n5904;
  assign n5906 = ~n5858 & ~n5905;
  assign n5907 = n5906 ^ n5867;
  assign n5908 = n5803 & ~n5905;
  assign n5909 = n5908 ^ n5805;
  assign n5910 = n5909 ^ n905;
  assign n5911 = n5796 & ~n5905;
  assign n5912 = n5911 ^ n5799;
  assign n5913 = n5912 ^ n1027;
  assign n5914 = n5755 ^ n2374;
  assign n5915 = ~n5905 & n5914;
  assign n5916 = n5915 ^ n5642;
  assign n5917 = n5916 ^ n2194;
  assign n5918 = n5752 ^ n2583;
  assign n5919 = ~n5905 & n5918;
  assign n5920 = n5919 ^ n5646;
  assign n5921 = n5920 ^ n2374;
  assign n5922 = n5711 & ~n5905;
  assign n5923 = n5922 ^ n5713;
  assign n5924 = n5923 ^ n3882;
  assign n5925 = n5705 & ~n5905;
  assign n5926 = n5925 ^ n5707;
  assign n5927 = n5926 ^ n4133;
  assign n5928 = ~x52 & ~x53;
  assign n5929 = ~n5625 & n5928;
  assign n5930 = ~x54 & n5929;
  assign n5931 = n5905 ^ x55;
  assign n5932 = x54 & n5625;
  assign n5933 = n5625 & ~n5928;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = n5934 ^ x54;
  assign n5936 = n5935 ^ n5934;
  assign n5937 = n5934 ^ n5905;
  assign n5938 = n5937 ^ n5934;
  assign n5939 = n5936 & ~n5938;
  assign n5940 = n5939 ^ n5934;
  assign n5941 = ~n5931 & n5940;
  assign n5942 = n5941 ^ n5934;
  assign n5943 = ~n5930 & ~n5942;
  assign n5944 = n5943 ^ n5363;
  assign n5945 = n5648 ^ n5625;
  assign n5946 = ~n5905 & ~n5945;
  assign n5947 = n5946 ^ n5625;
  assign n5948 = n5947 ^ x56;
  assign n5949 = n5948 ^ n5943;
  assign n5950 = n5944 & n5949;
  assign n5951 = n5950 ^ n5363;
  assign n5952 = n5951 ^ n5108;
  assign n5954 = n5652 ^ n5650;
  assign n5955 = n5954 ^ n5652;
  assign n5956 = n5654 ^ n5652;
  assign n5957 = n5956 ^ n5652;
  assign n5958 = ~n5955 & n5957;
  assign n5959 = n5958 ^ n5652;
  assign n5960 = n5625 & n5959;
  assign n5961 = n5960 ^ n5652;
  assign n5953 = ~x56 & ~n5625;
  assign n5962 = n5961 ^ n5953;
  assign n5963 = n5648 ^ n5363;
  assign n5964 = n5963 ^ n5961;
  assign n5965 = n5961 ^ n5905;
  assign n5966 = ~n5961 & n5965;
  assign n5967 = n5966 ^ n5961;
  assign n5968 = ~n5964 & ~n5967;
  assign n5969 = n5968 ^ n5966;
  assign n5970 = n5969 ^ n5961;
  assign n5971 = n5970 ^ n5905;
  assign n5972 = n5962 & n5971;
  assign n5973 = n5972 ^ n5953;
  assign n5974 = n5973 ^ x57;
  assign n5975 = n5974 ^ n5951;
  assign n5976 = n5952 & ~n5975;
  assign n5977 = n5976 ^ n5108;
  assign n5978 = n5977 ^ n4851;
  assign n5979 = n5664 & ~n5905;
  assign n5980 = n5979 ^ n5668;
  assign n5981 = n5980 ^ n5977;
  assign n5982 = n5978 & n5981;
  assign n5983 = n5982 ^ n4851;
  assign n5984 = n5983 ^ n4606;
  assign n5985 = n5672 & ~n5905;
  assign n5986 = n5985 ^ n5694;
  assign n5987 = n5986 ^ n5983;
  assign n5988 = n5984 & ~n5987;
  assign n5989 = n5988 ^ n4606;
  assign n5990 = n5989 ^ n4362;
  assign n5991 = n5698 & ~n5905;
  assign n5992 = n5991 ^ n5701;
  assign n5993 = n5992 ^ n5989;
  assign n5994 = n5990 & n5993;
  assign n5995 = n5994 ^ n4362;
  assign n5996 = n5995 ^ n5926;
  assign n5997 = n5927 & ~n5996;
  assign n5998 = n5997 ^ n4133;
  assign n5999 = n5998 ^ n5923;
  assign n6000 = ~n5924 & n5999;
  assign n6001 = n6000 ^ n3882;
  assign n6002 = n6001 ^ n3634;
  assign n6003 = n5717 & ~n5905;
  assign n6004 = n6003 ^ n5719;
  assign n6005 = n6004 ^ n6001;
  assign n6006 = ~n6002 & ~n6005;
  assign n6007 = n6006 ^ n3634;
  assign n6008 = n6007 ^ n3397;
  assign n6009 = ~n5723 & ~n5905;
  assign n6010 = n6009 ^ n5725;
  assign n6011 = n6010 ^ n6007;
  assign n6012 = ~n6008 & ~n6011;
  assign n6013 = n6012 ^ n3397;
  assign n6014 = n6013 ^ n3177;
  assign n6015 = ~n5729 & ~n5905;
  assign n6016 = n6015 ^ n5731;
  assign n6017 = n6016 ^ n6013;
  assign n6018 = n6014 & ~n6017;
  assign n6019 = n6018 ^ n3177;
  assign n6020 = n6019 ^ n2980;
  assign n6021 = n5735 & ~n5905;
  assign n6022 = n6021 ^ n5737;
  assign n6023 = n6022 ^ n6019;
  assign n6024 = n6020 & n6023;
  assign n6025 = n6024 ^ n2980;
  assign n6026 = n6025 ^ n2782;
  assign n6027 = n5741 & ~n5905;
  assign n6028 = n6027 ^ n5743;
  assign n6029 = n6028 ^ n6025;
  assign n6030 = n6026 & ~n6029;
  assign n6031 = n6030 ^ n2782;
  assign n6032 = n6031 ^ n2583;
  assign n6033 = n5747 & ~n5905;
  assign n6034 = n6033 ^ n5749;
  assign n6035 = n6034 ^ n6031;
  assign n6036 = n6032 & n6035;
  assign n6037 = n6036 ^ n2583;
  assign n6038 = n6037 ^ n5920;
  assign n6039 = n5921 & ~n6038;
  assign n6040 = n6039 ^ n2374;
  assign n6041 = n6040 ^ n5916;
  assign n6042 = n5917 & n6041;
  assign n6043 = n6042 ^ n2194;
  assign n6044 = n6043 ^ n2011;
  assign n6045 = ~n5759 & ~n5905;
  assign n6046 = n6045 ^ n5761;
  assign n6047 = n6046 ^ n6043;
  assign n6048 = ~n6044 & n6047;
  assign n6049 = n6048 ^ n2011;
  assign n6050 = n6049 ^ n1804;
  assign n6051 = ~n5765 & ~n5905;
  assign n6052 = n6051 ^ n5767;
  assign n6053 = n6052 ^ n6049;
  assign n6054 = n6050 & ~n6053;
  assign n6055 = n6054 ^ n1804;
  assign n6056 = n6055 ^ n1621;
  assign n6057 = n5771 & ~n5905;
  assign n6058 = n6057 ^ n5773;
  assign n6059 = n6058 ^ n6055;
  assign n6060 = n6056 & ~n6059;
  assign n6061 = n6060 ^ n1621;
  assign n6062 = n6061 ^ n1458;
  assign n6063 = n5777 & ~n5905;
  assign n6064 = n6063 ^ n5779;
  assign n6065 = n6064 ^ n6061;
  assign n6066 = n6062 & n6065;
  assign n6067 = n6066 ^ n1458;
  assign n6068 = n6067 ^ n1299;
  assign n6069 = n5783 & ~n5905;
  assign n6070 = n6069 ^ n5785;
  assign n6071 = n6070 ^ n6067;
  assign n6072 = n6068 & ~n6071;
  assign n6073 = n6072 ^ n1299;
  assign n6074 = n6073 ^ n1158;
  assign n6075 = n5789 & ~n5905;
  assign n6076 = n6075 ^ n5792;
  assign n6077 = n6076 ^ n6073;
  assign n6078 = n6074 & n6077;
  assign n6079 = n6078 ^ n1158;
  assign n6080 = n6079 ^ n5912;
  assign n6081 = n5913 & ~n6080;
  assign n6082 = n6081 ^ n1027;
  assign n6083 = n6082 ^ n5909;
  assign n6084 = n5910 & ~n6083;
  assign n6085 = n6084 ^ n905;
  assign n6086 = n6085 ^ n803;
  assign n6087 = n5808 ^ n905;
  assign n6088 = ~n5905 & n6087;
  assign n6089 = n6088 ^ n5638;
  assign n6090 = n6089 ^ n6085;
  assign n6091 = n6086 & ~n6090;
  assign n6092 = n6091 ^ n803;
  assign n6093 = n6092 ^ n707;
  assign n6094 = n5811 ^ n803;
  assign n6095 = ~n5905 & n6094;
  assign n6096 = n6095 ^ n5635;
  assign n6097 = n6096 ^ n6092;
  assign n6098 = ~n6093 & n6097;
  assign n6099 = n6098 ^ n707;
  assign n6100 = n6099 ^ n608;
  assign n6101 = ~n5815 & ~n5905;
  assign n6102 = n6101 ^ n5817;
  assign n6103 = n6102 ^ n6099;
  assign n6104 = ~n6100 & n6103;
  assign n6105 = n6104 ^ n608;
  assign n6106 = n6105 ^ n514;
  assign n6107 = ~n5821 & ~n5905;
  assign n6108 = n6107 ^ n5823;
  assign n6109 = n6108 ^ n6105;
  assign n6110 = n6106 & n6109;
  assign n6111 = n6110 ^ n514;
  assign n6112 = n6111 ^ n436;
  assign n6113 = n5827 & ~n5905;
  assign n6114 = n6113 ^ n5829;
  assign n6115 = n6114 ^ n6111;
  assign n6116 = n6112 & ~n6115;
  assign n6117 = n6116 ^ n436;
  assign n6118 = n6117 ^ n363;
  assign n6119 = n5833 & ~n5905;
  assign n6120 = n6119 ^ n5835;
  assign n6121 = n6120 ^ n6117;
  assign n6122 = n6118 & n6121;
  assign n6123 = n6122 ^ n363;
  assign n6124 = n6123 ^ n300;
  assign n6125 = n5838 ^ n363;
  assign n6126 = ~n5905 & n6125;
  assign n6127 = n6126 ^ n5632;
  assign n6128 = n6127 ^ n6123;
  assign n6129 = n6124 & ~n6128;
  assign n6130 = n6129 ^ n300;
  assign n6131 = n6130 ^ n243;
  assign n6132 = n5841 ^ n300;
  assign n6133 = ~n5905 & n6132;
  assign n6134 = n6133 ^ n5628;
  assign n6135 = n6134 ^ n6130;
  assign n6136 = n6131 & ~n6135;
  assign n6137 = n6136 ^ n243;
  assign n6138 = n6137 ^ n210;
  assign n6139 = n5845 & ~n5905;
  assign n6140 = n6139 ^ n5847;
  assign n6141 = n6140 ^ n6137;
  assign n6142 = n6138 & ~n6141;
  assign n6143 = n6142 ^ n210;
  assign n6144 = n6143 ^ n147;
  assign n6145 = n5851 & ~n5905;
  assign n6146 = n6145 ^ n5854;
  assign n6147 = n6146 ^ n6143;
  assign n6148 = ~n6144 & n6147;
  assign n6149 = n6148 ^ n147;
  assign n6150 = ~n5907 & n6149;
  assign n6151 = ~n132 & ~n6150;
  assign n6152 = n5907 & ~n6149;
  assign n6153 = ~n6151 & ~n6152;
  assign n6154 = n5871 & ~n5905;
  assign n6155 = n6154 ^ n5873;
  assign n6156 = ~n133 & n6155;
  assign n6157 = ~n6153 & ~n6156;
  assign n6158 = ~n133 & ~n5876;
  assign n6160 = n5873 & ~n5904;
  assign n6161 = n1292 & n6160;
  assign n6162 = n5870 & n6161;
  assign n6163 = ~n6158 & ~n6162;
  assign n6159 = ~n5904 & n6158;
  assign n6164 = n6163 ^ n6159;
  assign n6165 = n6164 ^ n6163;
  assign n6166 = n5873 ^ n5871;
  assign n6167 = n6166 ^ n5904;
  assign n6168 = ~n5870 & n6160;
  assign n6169 = n6168 ^ n5904;
  assign n6170 = n6169 ^ n5904;
  assign n6171 = n6170 ^ n5873;
  assign n6172 = n6167 & n6171;
  assign n6173 = n6172 ^ n6166;
  assign n6174 = n133 & ~n6173;
  assign n6175 = n6174 ^ n6163;
  assign n6176 = n6175 ^ n6163;
  assign n6177 = ~n6165 & ~n6176;
  assign n6178 = n6177 ^ n6163;
  assign n6179 = ~n5860 & ~n6178;
  assign n6180 = n6179 ^ n6163;
  assign n6181 = ~n6157 & ~n6180;
  assign n6182 = n6149 ^ n132;
  assign n6183 = ~n6181 & n6182;
  assign n6184 = n6183 ^ n5907;
  assign n6185 = ~n133 & ~n6184;
  assign n6186 = n6131 & ~n6181;
  assign n6187 = n6186 ^ n6134;
  assign n6188 = ~n210 & ~n6187;
  assign n6189 = n6138 & ~n6181;
  assign n6190 = n6189 ^ n6140;
  assign n6191 = n147 & ~n6190;
  assign n6192 = ~n6188 & ~n6191;
  assign n6193 = n6124 & ~n6181;
  assign n6194 = n6193 ^ n6127;
  assign n6195 = n6194 ^ n243;
  assign n6196 = n6112 & ~n6181;
  assign n6197 = n6196 ^ n6114;
  assign n6198 = ~n363 & ~n6197;
  assign n6199 = n6106 & ~n6181;
  assign n6200 = n6199 ^ n6108;
  assign n6201 = ~n436 & n6200;
  assign n6202 = ~n6198 & ~n6201;
  assign n6203 = n6074 & ~n6181;
  assign n6204 = n6203 ^ n6076;
  assign n6205 = n6204 ^ n1027;
  assign n6206 = n6068 & ~n6181;
  assign n6207 = n6206 ^ n6070;
  assign n6208 = n6207 ^ n1158;
  assign n6209 = n6062 & ~n6181;
  assign n6210 = n6209 ^ n6064;
  assign n6211 = n1299 & ~n6210;
  assign n6212 = n6211 ^ n6207;
  assign n6213 = n6208 & n6212;
  assign n6214 = n6213 ^ n6207;
  assign n6215 = n6214 ^ n6204;
  assign n6216 = n6215 ^ n6204;
  assign n6217 = ~n1158 & ~n6207;
  assign n6218 = ~n1299 & n6210;
  assign n6219 = ~n6217 & ~n6218;
  assign n6220 = n5984 & ~n6181;
  assign n6221 = n6220 ^ n5986;
  assign n6222 = n6221 ^ n4362;
  assign n6223 = n5978 & ~n6181;
  assign n6224 = n6223 ^ n5980;
  assign n6225 = n6224 ^ n4606;
  assign n6226 = n5928 ^ n5905;
  assign n6227 = ~n6181 & ~n6226;
  assign n6228 = n6227 ^ n5905;
  assign n6229 = n6228 ^ x54;
  assign n6230 = n6229 ^ n5625;
  assign n6231 = ~x50 & ~x51;
  assign n6232 = ~n5905 & n6231;
  assign n6233 = ~x52 & n6232;
  assign n6234 = n5905 & n6231;
  assign n6235 = ~x52 & n6234;
  assign n6236 = n6235 ^ n5905;
  assign n6237 = n6236 ^ n6181;
  assign n6238 = n6237 ^ x53;
  assign n6239 = n6238 ^ n6181;
  assign n6240 = n6239 ^ n6237;
  assign n6241 = ~x52 & ~n6181;
  assign n6242 = n6241 ^ n6237;
  assign n6243 = ~n6240 & ~n6242;
  assign n6244 = n6243 ^ n6238;
  assign n6245 = ~n6233 & ~n6244;
  assign n6246 = n6245 ^ n6229;
  assign n6247 = ~n6230 & n6246;
  assign n6248 = n6247 ^ n5625;
  assign n6249 = n6248 ^ n5363;
  assign n6251 = n5932 ^ n5930;
  assign n6252 = n6251 ^ n5932;
  assign n6253 = n5934 ^ n5932;
  assign n6254 = n6253 ^ n5932;
  assign n6255 = ~n6252 & n6254;
  assign n6256 = n6255 ^ n5932;
  assign n6257 = n5905 & n6256;
  assign n6258 = n6257 ^ n5932;
  assign n6250 = ~x54 & ~n5905;
  assign n6259 = n6258 ^ n6250;
  assign n6260 = n5928 ^ n5625;
  assign n6261 = n6260 ^ n6258;
  assign n6262 = n6258 ^ n6181;
  assign n6263 = ~n6258 & n6262;
  assign n6264 = n6263 ^ n6258;
  assign n6265 = ~n6261 & ~n6264;
  assign n6266 = n6265 ^ n6263;
  assign n6267 = n6266 ^ n6258;
  assign n6268 = n6267 ^ n6181;
  assign n6269 = n6259 & n6268;
  assign n6270 = n6269 ^ n6250;
  assign n6271 = n6270 ^ x55;
  assign n6272 = n6271 ^ n6248;
  assign n6273 = n6249 & ~n6272;
  assign n6274 = n6273 ^ n5363;
  assign n6275 = n6274 ^ n5108;
  assign n6276 = n5944 & ~n6181;
  assign n6277 = n6276 ^ n5948;
  assign n6278 = n6277 ^ n6274;
  assign n6279 = n6275 & n6278;
  assign n6280 = n6279 ^ n5108;
  assign n6281 = n6280 ^ n4851;
  assign n6282 = n5952 & ~n6181;
  assign n6283 = n6282 ^ n5974;
  assign n6284 = n6283 ^ n6280;
  assign n6285 = n6281 & ~n6284;
  assign n6286 = n6285 ^ n4851;
  assign n6287 = n6286 ^ n6224;
  assign n6288 = ~n6225 & n6287;
  assign n6289 = n6288 ^ n4606;
  assign n6290 = n6289 ^ n6221;
  assign n6291 = n6222 & ~n6290;
  assign n6292 = n6291 ^ n4362;
  assign n6293 = n6292 ^ n4133;
  assign n6294 = n5990 & ~n6181;
  assign n6295 = n6294 ^ n5992;
  assign n6296 = n6295 ^ n6292;
  assign n6297 = n6293 & n6296;
  assign n6298 = n6297 ^ n4133;
  assign n6299 = n6298 ^ n3882;
  assign n6300 = n5995 ^ n4133;
  assign n6301 = ~n6181 & n6300;
  assign n6302 = n6301 ^ n5926;
  assign n6303 = n6302 ^ n6298;
  assign n6304 = n6299 & ~n6303;
  assign n6305 = n6304 ^ n3882;
  assign n6306 = n6305 ^ n3634;
  assign n6307 = n5998 ^ n3882;
  assign n6308 = ~n6181 & n6307;
  assign n6309 = n6308 ^ n5923;
  assign n6310 = n6309 ^ n6305;
  assign n6311 = ~n6306 & n6310;
  assign n6312 = n6311 ^ n3634;
  assign n6313 = n6312 ^ n3397;
  assign n6314 = ~n6002 & ~n6181;
  assign n6315 = n6314 ^ n6004;
  assign n6316 = n6315 ^ n6312;
  assign n6317 = ~n6313 & n6316;
  assign n6318 = n6317 ^ n3397;
  assign n6319 = n6318 ^ n3177;
  assign n6320 = ~n6008 & ~n6181;
  assign n6321 = n6320 ^ n6010;
  assign n6322 = n6321 ^ n6318;
  assign n6323 = n6319 & n6322;
  assign n6324 = n6323 ^ n3177;
  assign n6325 = n6324 ^ n2980;
  assign n6326 = n6014 & ~n6181;
  assign n6327 = n6326 ^ n6016;
  assign n6328 = n6327 ^ n6324;
  assign n6329 = n6325 & ~n6328;
  assign n6330 = n6329 ^ n2980;
  assign n6331 = n6330 ^ n2782;
  assign n6332 = n6020 & ~n6181;
  assign n6333 = n6332 ^ n6022;
  assign n6334 = n6333 ^ n6330;
  assign n6335 = n6331 & n6334;
  assign n6336 = n6335 ^ n2782;
  assign n6337 = n6336 ^ n2583;
  assign n6338 = n6026 & ~n6181;
  assign n6339 = n6338 ^ n6028;
  assign n6340 = n6339 ^ n6336;
  assign n6341 = n6337 & ~n6340;
  assign n6342 = n6341 ^ n2583;
  assign n6343 = n6342 ^ n2374;
  assign n6344 = n6032 & ~n6181;
  assign n6345 = n6344 ^ n6034;
  assign n6346 = n6345 ^ n6342;
  assign n6347 = n6343 & n6346;
  assign n6348 = n6347 ^ n2374;
  assign n6349 = n6348 ^ n2194;
  assign n6350 = n6037 ^ n2374;
  assign n6351 = ~n6181 & n6350;
  assign n6352 = n6351 ^ n5920;
  assign n6353 = n6352 ^ n6348;
  assign n6354 = ~n6349 & ~n6353;
  assign n6355 = n6354 ^ n2194;
  assign n6356 = n6355 ^ n2011;
  assign n6357 = n6040 ^ n2194;
  assign n6358 = ~n6181 & ~n6357;
  assign n6359 = n6358 ^ n5916;
  assign n6360 = n6359 ^ n6355;
  assign n6361 = ~n6356 & ~n6360;
  assign n6362 = n6361 ^ n2011;
  assign n6363 = n6362 ^ n1804;
  assign n6364 = ~n6044 & ~n6181;
  assign n6365 = n6364 ^ n6046;
  assign n6366 = n6365 ^ n6362;
  assign n6367 = n6363 & ~n6366;
  assign n6368 = n6367 ^ n1804;
  assign n6369 = n6368 ^ n1621;
  assign n6370 = n6050 & ~n6181;
  assign n6371 = n6370 ^ n6052;
  assign n6372 = n6371 ^ n6368;
  assign n6373 = n6369 & ~n6372;
  assign n6374 = n6373 ^ n1621;
  assign n6375 = n6374 ^ n1458;
  assign n6376 = n6056 & ~n6181;
  assign n6377 = n6376 ^ n6058;
  assign n6378 = n6377 ^ n6374;
  assign n6379 = n6375 & ~n6378;
  assign n6380 = n6379 ^ n1458;
  assign n6381 = n6219 & n6380;
  assign n6382 = n6381 ^ n6204;
  assign n6383 = n6382 ^ n6204;
  assign n6384 = ~n6216 & ~n6383;
  assign n6385 = n6384 ^ n6204;
  assign n6386 = ~n6205 & ~n6385;
  assign n6387 = n6386 ^ n1027;
  assign n6388 = n6387 ^ n905;
  assign n6389 = n6079 ^ n1027;
  assign n6390 = ~n6181 & n6389;
  assign n6391 = n6390 ^ n5912;
  assign n6392 = n6391 ^ n6387;
  assign n6393 = n6388 & ~n6392;
  assign n6394 = n6393 ^ n905;
  assign n6395 = n6394 ^ n803;
  assign n6396 = n6082 ^ n905;
  assign n6397 = ~n6181 & n6396;
  assign n6398 = n6397 ^ n5909;
  assign n6399 = n6398 ^ n6394;
  assign n6400 = n6395 & ~n6399;
  assign n6401 = n6400 ^ n803;
  assign n6402 = n6401 ^ n707;
  assign n6403 = n6086 & ~n6181;
  assign n6404 = n6403 ^ n6089;
  assign n6405 = n6404 ^ n6401;
  assign n6406 = ~n6402 & ~n6405;
  assign n6407 = n6406 ^ n707;
  assign n6408 = n6407 ^ n608;
  assign n6409 = ~n6093 & ~n6181;
  assign n6410 = n6409 ^ n6096;
  assign n6411 = n6410 ^ n6407;
  assign n6412 = ~n6408 & ~n6411;
  assign n6413 = n6412 ^ n608;
  assign n6414 = n6413 ^ n514;
  assign n6415 = ~n6100 & ~n6181;
  assign n6416 = n6415 ^ n6102;
  assign n6417 = n6416 ^ n6413;
  assign n6418 = n6414 & ~n6417;
  assign n6419 = n6418 ^ n514;
  assign n6420 = n6202 & n6419;
  assign n6421 = n6197 ^ n363;
  assign n6422 = n436 & ~n6200;
  assign n6423 = n6422 ^ n6197;
  assign n6424 = n6421 & ~n6423;
  assign n6425 = n6424 ^ n363;
  assign n6426 = ~n6420 & ~n6425;
  assign n6427 = n6426 ^ n300;
  assign n6428 = n6118 & ~n6181;
  assign n6429 = n6428 ^ n6120;
  assign n6430 = n6429 ^ n6426;
  assign n6431 = ~n6427 & ~n6430;
  assign n6432 = n6431 ^ n300;
  assign n6433 = n6432 ^ n6194;
  assign n6434 = n6195 & ~n6433;
  assign n6435 = n6434 ^ n243;
  assign n6436 = n6192 & n6435;
  assign n6437 = n6190 ^ n147;
  assign n6438 = n210 & n6187;
  assign n6439 = n6438 ^ n6190;
  assign n6440 = ~n6437 & ~n6439;
  assign n6441 = n6440 ^ n147;
  assign n6442 = ~n6436 & n6441;
  assign n6443 = n6442 ^ n132;
  assign n6444 = ~n6144 & ~n6181;
  assign n6445 = n6444 ^ n6146;
  assign n6446 = n6445 ^ n6442;
  assign n6447 = n6443 & ~n6446;
  assign n6448 = n6447 ^ n132;
  assign n6449 = ~n6185 & ~n6448;
  assign n6450 = ~n132 & n6149;
  assign n6451 = ~n5907 & ~n6155;
  assign n6452 = n6450 & n6451;
  assign n6453 = n6150 & n6180;
  assign n6454 = n6155 & ~n6453;
  assign n6455 = n132 & n6180;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = ~n132 & n5907;
  assign n6458 = n6155 & ~n6457;
  assign n6459 = ~n6149 & ~n6458;
  assign n6460 = n6149 ^ n5907;
  assign n6461 = n6460 ^ n6149;
  assign n6462 = n6155 & n6180;
  assign n6463 = n6462 ^ n6149;
  assign n6464 = ~n6461 & n6463;
  assign n6465 = n6464 ^ n6149;
  assign n6466 = n132 & n6465;
  assign n6467 = ~n6459 & ~n6466;
  assign n6468 = ~n6456 & n6467;
  assign n6469 = n6468 ^ n133;
  assign n6470 = n6469 ^ n6468;
  assign n6471 = ~n6153 & n6462;
  assign n6472 = n132 & ~n6155;
  assign n6473 = ~n6152 & n6472;
  assign n6474 = ~n6471 & ~n6473;
  assign n6475 = n6474 ^ n6468;
  assign n6476 = ~n6470 & n6475;
  assign n6477 = n6476 ^ n6468;
  assign n6478 = ~n6452 & n6477;
  assign n6479 = ~n6449 & n6478;
  assign n6480 = n6435 ^ n210;
  assign n6481 = n6435 ^ n6187;
  assign n6482 = n6480 & ~n6481;
  assign n6483 = n6482 ^ n210;
  assign n6484 = n6483 ^ n147;
  assign n6485 = ~n6479 & ~n6484;
  assign n6486 = n6485 ^ n6190;
  assign n6487 = ~n6479 & n6480;
  assign n6488 = n6487 ^ n6187;
  assign n6489 = n6488 ^ n147;
  assign n6490 = n6414 & ~n6479;
  assign n6491 = n6490 ^ n6416;
  assign n6492 = n6491 ^ n436;
  assign n6493 = ~n6408 & ~n6479;
  assign n6494 = n6493 ^ n6410;
  assign n6495 = n6494 ^ n514;
  assign n6496 = ~n6402 & ~n6479;
  assign n6497 = n6496 ^ n6404;
  assign n6498 = n608 & n6497;
  assign n6499 = n6498 ^ n6494;
  assign n6500 = ~n6495 & ~n6499;
  assign n6501 = n6500 ^ n6494;
  assign n6502 = n6501 ^ n6491;
  assign n6503 = n6502 ^ n6491;
  assign n6504 = ~n608 & ~n6497;
  assign n6505 = ~n514 & n6494;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = n6369 & ~n6479;
  assign n6508 = n6507 ^ n6371;
  assign n6509 = n6508 ^ n1458;
  assign n6510 = n6363 & ~n6479;
  assign n6511 = n6510 ^ n6365;
  assign n6512 = n6511 ^ n1621;
  assign n6513 = n6299 & ~n6479;
  assign n6514 = n6513 ^ n6302;
  assign n6515 = n6514 ^ n3634;
  assign n6516 = n6293 & ~n6479;
  assign n6517 = n6516 ^ n6295;
  assign n6518 = n6517 ^ n3882;
  assign n6519 = x50 & ~n6479;
  assign n6520 = ~x51 & n6519;
  assign n6521 = ~x48 & ~x49;
  assign n6522 = ~n6181 & n6521;
  assign n6523 = ~x50 & n6522;
  assign n6524 = ~n6520 & ~n6523;
  assign n6525 = n6181 & ~n6521;
  assign n6526 = x50 & n6181;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = n6479 ^ x51;
  assign n6529 = n6527 & n6528;
  assign n6530 = n6524 & ~n6529;
  assign n6531 = n6530 ^ n5905;
  assign n6532 = n6231 ^ n6181;
  assign n6533 = ~n6479 & ~n6532;
  assign n6534 = n6533 ^ n6181;
  assign n6535 = n6534 ^ x52;
  assign n6536 = n6535 ^ n6530;
  assign n6537 = n6531 & n6536;
  assign n6538 = n6537 ^ n5905;
  assign n6539 = n6538 ^ n5625;
  assign n6540 = n6181 ^ n5905;
  assign n6541 = n6540 ^ n6181;
  assign n6542 = n6541 ^ n6540;
  assign n6543 = n6540 ^ n6231;
  assign n6544 = n6542 & n6543;
  assign n6545 = n6544 ^ n6540;
  assign n6546 = ~x52 & n6545;
  assign n6547 = n6546 ^ n6540;
  assign n6548 = n6547 ^ n6241;
  assign n6549 = n6231 ^ n5905;
  assign n6550 = n6549 ^ n6547;
  assign n6551 = n6547 ^ n6479;
  assign n6552 = ~n6547 & n6551;
  assign n6553 = n6552 ^ n6547;
  assign n6554 = ~n6550 & ~n6553;
  assign n6555 = n6554 ^ n6552;
  assign n6556 = n6555 ^ n6547;
  assign n6557 = n6556 ^ n6479;
  assign n6558 = n6548 & n6557;
  assign n6559 = n6558 ^ n6241;
  assign n6560 = n6559 ^ x53;
  assign n6561 = n6560 ^ n6538;
  assign n6562 = n6539 & ~n6561;
  assign n6563 = n6562 ^ n5625;
  assign n6564 = n6563 ^ n5363;
  assign n6565 = n6245 ^ n5625;
  assign n6566 = ~n6479 & n6565;
  assign n6567 = n6566 ^ n6229;
  assign n6568 = n6567 ^ n6563;
  assign n6569 = n6564 & n6568;
  assign n6570 = n6569 ^ n5363;
  assign n6571 = n6570 ^ n5108;
  assign n6572 = n6249 & ~n6479;
  assign n6573 = n6572 ^ n6271;
  assign n6574 = n6573 ^ n6570;
  assign n6575 = n6571 & ~n6574;
  assign n6576 = n6575 ^ n5108;
  assign n6577 = n6576 ^ n4851;
  assign n6578 = n6275 & ~n6479;
  assign n6579 = n6578 ^ n6277;
  assign n6580 = n6579 ^ n6576;
  assign n6581 = n6577 & n6580;
  assign n6582 = n6581 ^ n4851;
  assign n6583 = n6582 ^ n4606;
  assign n6584 = n6281 & ~n6479;
  assign n6585 = n6584 ^ n6283;
  assign n6586 = n6585 ^ n6582;
  assign n6587 = n6583 & ~n6586;
  assign n6588 = n6587 ^ n4606;
  assign n6589 = n6588 ^ n4362;
  assign n6590 = n6286 ^ n4606;
  assign n6591 = ~n6479 & n6590;
  assign n6592 = n6591 ^ n6224;
  assign n6593 = n6592 ^ n6588;
  assign n6594 = n6589 & n6593;
  assign n6595 = n6594 ^ n4362;
  assign n6596 = n6595 ^ n4133;
  assign n6597 = n6289 ^ n4362;
  assign n6598 = ~n6479 & n6597;
  assign n6599 = n6598 ^ n6221;
  assign n6600 = n6599 ^ n6595;
  assign n6601 = n6596 & ~n6600;
  assign n6602 = n6601 ^ n4133;
  assign n6603 = n6602 ^ n6517;
  assign n6604 = ~n6518 & n6603;
  assign n6605 = n6604 ^ n3882;
  assign n6606 = n6605 ^ n6514;
  assign n6607 = ~n6515 & ~n6606;
  assign n6608 = n6607 ^ n3634;
  assign n6609 = n6608 ^ n3397;
  assign n6610 = ~n6306 & ~n6479;
  assign n6611 = n6610 ^ n6309;
  assign n6612 = n6611 ^ n6608;
  assign n6613 = ~n6609 & ~n6612;
  assign n6614 = n6613 ^ n3397;
  assign n6615 = n6614 ^ n3177;
  assign n6616 = ~n6313 & ~n6479;
  assign n6617 = n6616 ^ n6315;
  assign n6618 = n6617 ^ n6614;
  assign n6619 = n6615 & ~n6618;
  assign n6620 = n6619 ^ n3177;
  assign n6621 = n6620 ^ n2980;
  assign n6622 = n6319 & ~n6479;
  assign n6623 = n6622 ^ n6321;
  assign n6624 = n6623 ^ n6620;
  assign n6625 = n6621 & n6624;
  assign n6626 = n6625 ^ n2980;
  assign n6627 = n6626 ^ n2782;
  assign n6628 = n6325 & ~n6479;
  assign n6629 = n6628 ^ n6327;
  assign n6630 = n6629 ^ n6626;
  assign n6631 = n6627 & ~n6630;
  assign n6632 = n6631 ^ n2782;
  assign n6633 = n6632 ^ n2583;
  assign n6634 = n6331 & ~n6479;
  assign n6635 = n6634 ^ n6333;
  assign n6636 = n6635 ^ n6632;
  assign n6637 = n6633 & n6636;
  assign n6638 = n6637 ^ n2583;
  assign n6639 = n6638 ^ n2374;
  assign n6640 = n6337 & ~n6479;
  assign n6641 = n6640 ^ n6339;
  assign n6642 = n6641 ^ n6638;
  assign n6643 = n6639 & ~n6642;
  assign n6644 = n6643 ^ n2374;
  assign n6645 = n6644 ^ n2194;
  assign n6646 = n6343 & ~n6479;
  assign n6647 = n6646 ^ n6345;
  assign n6648 = n6647 ^ n6644;
  assign n6649 = ~n6645 & n6648;
  assign n6650 = n6649 ^ n2194;
  assign n6651 = n6650 ^ n2011;
  assign n6652 = ~n6349 & ~n6479;
  assign n6653 = n6652 ^ n6352;
  assign n6654 = n6653 ^ n6650;
  assign n6655 = ~n6651 & n6654;
  assign n6656 = n6655 ^ n2011;
  assign n6657 = n6656 ^ n1804;
  assign n6658 = ~n6356 & ~n6479;
  assign n6659 = n6658 ^ n6359;
  assign n6660 = n6659 ^ n6656;
  assign n6661 = n6657 & n6660;
  assign n6662 = n6661 ^ n1804;
  assign n6663 = n6662 ^ n6511;
  assign n6664 = n6512 & ~n6663;
  assign n6665 = n6664 ^ n1621;
  assign n6666 = n6665 ^ n6508;
  assign n6667 = n6509 & ~n6666;
  assign n6668 = n6667 ^ n1458;
  assign n6669 = n6668 ^ n1299;
  assign n6670 = n6375 & ~n6479;
  assign n6671 = n6670 ^ n6377;
  assign n6672 = n6671 ^ n6668;
  assign n6673 = n6669 & ~n6672;
  assign n6674 = n6673 ^ n1299;
  assign n6675 = n6674 ^ n1158;
  assign n6676 = n6380 ^ n1299;
  assign n6677 = ~n6479 & n6676;
  assign n6678 = n6677 ^ n6210;
  assign n6679 = n6678 ^ n6674;
  assign n6680 = n6675 & n6679;
  assign n6681 = n6680 ^ n1158;
  assign n6682 = n6681 ^ n1027;
  assign n6683 = n6210 ^ n1299;
  assign n6684 = n6380 ^ n6210;
  assign n6685 = ~n6683 & n6684;
  assign n6686 = n6685 ^ n1299;
  assign n6687 = n6686 ^ n1158;
  assign n6688 = ~n6479 & n6687;
  assign n6689 = n6688 ^ n6207;
  assign n6690 = n6689 ^ n6681;
  assign n6691 = n6682 & ~n6690;
  assign n6692 = n6691 ^ n1027;
  assign n6693 = n6692 ^ n905;
  assign n6694 = n6686 ^ n6207;
  assign n6695 = n6208 & ~n6694;
  assign n6696 = n6695 ^ n1158;
  assign n6697 = n6696 ^ n1027;
  assign n6698 = ~n6479 & n6697;
  assign n6699 = n6698 ^ n6204;
  assign n6700 = n6699 ^ n6692;
  assign n6701 = n6693 & n6700;
  assign n6702 = n6701 ^ n905;
  assign n6703 = n6702 ^ n803;
  assign n6704 = n6388 & ~n6479;
  assign n6705 = n6704 ^ n6391;
  assign n6706 = n6705 ^ n6702;
  assign n6707 = n6703 & ~n6706;
  assign n6708 = n6707 ^ n803;
  assign n6709 = n6708 ^ n707;
  assign n6710 = n6395 & ~n6479;
  assign n6711 = n6710 ^ n6398;
  assign n6712 = n6711 ^ n6708;
  assign n6713 = ~n6709 & ~n6712;
  assign n6714 = n6713 ^ n707;
  assign n6715 = n6506 & ~n6714;
  assign n6716 = n6715 ^ n6491;
  assign n6717 = n6716 ^ n6491;
  assign n6718 = n6503 & ~n6717;
  assign n6719 = n6718 ^ n6491;
  assign n6720 = n6492 & n6719;
  assign n6721 = n6720 ^ n436;
  assign n6722 = n6721 ^ n363;
  assign n6723 = n6419 ^ n436;
  assign n6724 = ~n6479 & n6723;
  assign n6725 = n6724 ^ n6200;
  assign n6726 = n6725 ^ n6721;
  assign n6727 = n6722 & n6726;
  assign n6728 = n6727 ^ n363;
  assign n6729 = n6728 ^ n300;
  assign n6730 = n6419 ^ n6200;
  assign n6731 = n6723 & n6730;
  assign n6732 = n6731 ^ n436;
  assign n6733 = n6732 ^ n363;
  assign n6734 = ~n6479 & n6733;
  assign n6735 = n6734 ^ n6197;
  assign n6736 = n6735 ^ n6728;
  assign n6737 = n6729 & ~n6736;
  assign n6738 = n6737 ^ n300;
  assign n6739 = n6738 ^ n243;
  assign n6740 = ~n6427 & ~n6479;
  assign n6741 = n6740 ^ n6429;
  assign n6742 = n6741 ^ n6738;
  assign n6743 = n6739 & n6742;
  assign n6744 = n6743 ^ n243;
  assign n6745 = n6744 ^ n210;
  assign n6746 = n6432 ^ n243;
  assign n6747 = ~n6479 & n6746;
  assign n6748 = n6747 ^ n6194;
  assign n6749 = n6748 ^ n6744;
  assign n6750 = n6745 & ~n6749;
  assign n6751 = n6750 ^ n210;
  assign n6752 = n6751 ^ n6488;
  assign n6753 = ~n6489 & ~n6752;
  assign n6754 = n6753 ^ n147;
  assign n6755 = n6486 & ~n6754;
  assign n6756 = ~n6486 & n6754;
  assign n6757 = ~n132 & ~n6756;
  assign n6758 = ~n6755 & ~n6757;
  assign n6759 = n6443 & ~n6479;
  assign n6760 = n6759 ^ n6445;
  assign n6761 = ~n133 & n6760;
  assign n6762 = ~n6758 & ~n6761;
  assign n6776 = ~n133 & ~n6448;
  assign n6777 = n6442 & n6445;
  assign n6778 = ~n6152 & n6155;
  assign n6779 = n6151 & n6778;
  assign n6780 = ~n5907 & n6155;
  assign n6781 = ~n6180 & n6780;
  assign n6782 = n1292 & ~n6781;
  assign n6783 = ~n6779 & n6782;
  assign n6784 = n6155 ^ n6152;
  assign n6785 = n6784 ^ n6152;
  assign n6786 = n6453 ^ n6152;
  assign n6787 = ~n6785 & n6786;
  assign n6788 = n6787 ^ n6152;
  assign n6789 = n132 & n6788;
  assign n6790 = n6783 & ~n6789;
  assign n6791 = n6777 & n6790;
  assign n6792 = ~n6776 & ~n6791;
  assign n6763 = n6445 ^ n6443;
  assign n6764 = n6763 ^ n6478;
  assign n6765 = n6478 ^ n6442;
  assign n6766 = n6478 ^ n6445;
  assign n6767 = ~n6478 & ~n6766;
  assign n6768 = n6767 ^ n6478;
  assign n6769 = n6765 & ~n6768;
  assign n6770 = n6769 ^ n6767;
  assign n6771 = n6770 ^ n6478;
  assign n6772 = n6771 ^ n6445;
  assign n6773 = n6764 & ~n6772;
  assign n6774 = n6773 ^ n6763;
  assign n6775 = n133 & ~n6774;
  assign n6793 = n6792 ^ n6775;
  assign n6794 = n6793 ^ n6792;
  assign n6795 = ~n6478 & n6776;
  assign n6796 = n6795 ^ n6792;
  assign n6797 = n6796 ^ n6792;
  assign n6798 = ~n6794 & ~n6797;
  assign n6799 = n6798 ^ n6792;
  assign n6800 = ~n6184 & ~n6799;
  assign n6801 = n6800 ^ n6792;
  assign n6802 = ~n6762 & ~n6801;
  assign n6803 = n6754 & n6802;
  assign n6804 = n6722 & ~n6802;
  assign n6805 = n6804 ^ n6725;
  assign n6806 = n6805 ^ n300;
  assign n6807 = n6497 ^ n608;
  assign n6808 = n6714 ^ n6497;
  assign n6809 = n6807 & n6808;
  assign n6810 = n6809 ^ n608;
  assign n6811 = n6810 ^ n6494;
  assign n6812 = ~n6495 & n6811;
  assign n6813 = n6812 ^ n514;
  assign n6814 = n6813 ^ n436;
  assign n6815 = ~n6802 & n6814;
  assign n6816 = n6815 ^ n6491;
  assign n6817 = n6816 ^ n363;
  assign n6818 = n6657 & ~n6802;
  assign n6819 = n6818 ^ n6659;
  assign n6820 = n6819 ^ n1621;
  assign n6821 = ~n6651 & ~n6802;
  assign n6822 = n6821 ^ n6653;
  assign n6823 = n6822 ^ n1804;
  assign n6824 = ~n6645 & ~n6802;
  assign n6825 = n6824 ^ n6647;
  assign n6826 = n2011 & ~n6825;
  assign n6827 = n6826 ^ n6822;
  assign n6828 = n6823 & n6827;
  assign n6829 = n6828 ^ n6822;
  assign n6830 = n6829 ^ n6819;
  assign n6831 = n6830 ^ n6819;
  assign n6832 = ~n1804 & ~n6822;
  assign n6833 = ~n2011 & n6825;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = n6627 & ~n6802;
  assign n6836 = n6835 ^ n6629;
  assign n6837 = n6836 ^ n2583;
  assign n6838 = n6621 & ~n6802;
  assign n6839 = n6838 ^ n6623;
  assign n6840 = n6839 ^ n2782;
  assign n6841 = n6615 & ~n6802;
  assign n6842 = n6841 ^ n6617;
  assign n6843 = ~n2980 & ~n6842;
  assign n6844 = n6843 ^ n6839;
  assign n6845 = ~n6840 & n6844;
  assign n6846 = n6845 ^ n6839;
  assign n6847 = n6846 ^ n6836;
  assign n6848 = n6847 ^ n6836;
  assign n6849 = n2980 & n6842;
  assign n6850 = n2782 & ~n6839;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = n6583 & ~n6802;
  assign n6853 = n6852 ^ n6585;
  assign n6854 = n6853 ^ n4362;
  assign n6855 = n6577 & ~n6802;
  assign n6856 = n6855 ^ n6579;
  assign n6857 = n6856 ^ n4606;
  assign n6858 = n6521 ^ n6479;
  assign n6859 = ~n6802 & ~n6858;
  assign n6860 = n6859 ^ n6479;
  assign n6861 = ~x50 & n6860;
  assign n6862 = ~x46 & ~x47;
  assign n6863 = ~n6479 & n6862;
  assign n6864 = ~x48 & n6863;
  assign n6865 = ~x48 & n6862;
  assign n6866 = ~x49 & x50;
  assign n6867 = n6865 & n6866;
  assign n6868 = ~n6519 & ~n6867;
  assign n6869 = ~n6864 & n6868;
  assign n6870 = n6802 ^ x50;
  assign n6871 = n6870 ^ x49;
  assign n6872 = x49 & ~n6802;
  assign n6873 = n6865 & n6872;
  assign n6874 = n6873 ^ n6870;
  assign n6875 = n6870 & ~n6874;
  assign n6876 = n6875 ^ n6870;
  assign n6877 = ~n6871 & n6876;
  assign n6878 = n6877 ^ n6875;
  assign n6879 = n6878 ^ n6870;
  assign n6880 = n6879 ^ n6873;
  assign n6881 = n6869 & ~n6880;
  assign n6882 = ~n6861 & n6881;
  assign n6883 = ~n6521 & ~n6802;
  assign n6884 = n6479 & ~n6862;
  assign n6885 = x48 & n6479;
  assign n6886 = ~n6884 & ~n6885;
  assign n6887 = x49 & ~n6886;
  assign n6888 = ~x50 & ~n6887;
  assign n6889 = n6883 & n6888;
  assign n6890 = x49 & ~n6864;
  assign n6891 = n6479 ^ x50;
  assign n6892 = n6479 & ~n6865;
  assign n6893 = n6891 & n6892;
  assign n6894 = n6893 ^ n6891;
  assign n6895 = ~n6890 & n6894;
  assign n6896 = n6802 & n6895;
  assign n6897 = ~n6479 & n6867;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = ~n6889 & n6898;
  assign n6900 = n6181 & n6899;
  assign n6901 = ~n6882 & ~n6900;
  assign n6902 = n6901 ^ n5905;
  assign n6904 = ~n6523 & n6527;
  assign n6905 = n6904 ^ n6526;
  assign n6906 = n6479 & n6905;
  assign n6907 = n6906 ^ n6526;
  assign n6903 = ~x50 & ~n6479;
  assign n6908 = n6907 ^ n6903;
  assign n6909 = n6521 ^ n6181;
  assign n6910 = n6909 ^ n6907;
  assign n6911 = n6907 ^ n6802;
  assign n6912 = ~n6907 & n6911;
  assign n6913 = n6912 ^ n6907;
  assign n6914 = ~n6910 & ~n6913;
  assign n6915 = n6914 ^ n6912;
  assign n6916 = n6915 ^ n6907;
  assign n6917 = n6916 ^ n6802;
  assign n6918 = n6908 & n6917;
  assign n6919 = n6918 ^ n6903;
  assign n6920 = n6919 ^ x51;
  assign n6921 = n6920 ^ n6901;
  assign n6922 = ~n6902 & n6921;
  assign n6923 = n6922 ^ n5905;
  assign n6924 = n6923 ^ n5625;
  assign n6925 = n6531 & ~n6802;
  assign n6926 = n6925 ^ n6535;
  assign n6927 = n6926 ^ n6923;
  assign n6928 = n6924 & n6927;
  assign n6929 = n6928 ^ n5625;
  assign n6930 = n6929 ^ n5363;
  assign n6931 = n6539 & ~n6802;
  assign n6932 = n6931 ^ n6560;
  assign n6933 = n6932 ^ n6929;
  assign n6934 = n6930 & ~n6933;
  assign n6935 = n6934 ^ n5363;
  assign n6936 = n6935 ^ n5108;
  assign n6937 = n6564 & ~n6802;
  assign n6938 = n6937 ^ n6567;
  assign n6939 = n6938 ^ n6935;
  assign n6940 = n6936 & n6939;
  assign n6941 = n6940 ^ n5108;
  assign n6942 = n6941 ^ n4851;
  assign n6943 = n6571 & ~n6802;
  assign n6944 = n6943 ^ n6573;
  assign n6945 = n6944 ^ n6941;
  assign n6946 = n6942 & ~n6945;
  assign n6947 = n6946 ^ n4851;
  assign n6948 = n6947 ^ n6856;
  assign n6949 = ~n6857 & n6948;
  assign n6950 = n6949 ^ n4606;
  assign n6951 = n6950 ^ n6853;
  assign n6952 = n6854 & ~n6951;
  assign n6953 = n6952 ^ n4362;
  assign n6954 = n6953 ^ n4133;
  assign n6955 = n6589 & ~n6802;
  assign n6956 = n6955 ^ n6592;
  assign n6957 = n6956 ^ n6953;
  assign n6958 = n6954 & n6957;
  assign n6959 = n6958 ^ n4133;
  assign n6960 = n6959 ^ n3882;
  assign n6961 = n6596 & ~n6802;
  assign n6962 = n6961 ^ n6599;
  assign n6963 = n6962 ^ n6959;
  assign n6964 = n6960 & ~n6963;
  assign n6965 = n6964 ^ n3882;
  assign n6966 = n6965 ^ n3634;
  assign n6967 = n6602 ^ n3882;
  assign n6968 = ~n6802 & n6967;
  assign n6969 = n6968 ^ n6517;
  assign n6970 = n6969 ^ n6965;
  assign n6971 = ~n6966 & n6970;
  assign n6972 = n6971 ^ n3634;
  assign n6973 = n6972 ^ n3397;
  assign n6974 = n6605 ^ n3634;
  assign n6975 = ~n6802 & ~n6974;
  assign n6976 = n6975 ^ n6514;
  assign n6977 = n6976 ^ n6972;
  assign n6978 = ~n6973 & n6977;
  assign n6979 = n6978 ^ n3397;
  assign n6980 = n6979 ^ n3177;
  assign n6981 = ~n6609 & ~n6802;
  assign n6982 = n6981 ^ n6611;
  assign n6983 = n6982 ^ n6979;
  assign n6984 = n6980 & n6983;
  assign n6985 = n6984 ^ n3177;
  assign n6986 = n6851 & ~n6985;
  assign n6987 = n6986 ^ n6836;
  assign n6988 = n6987 ^ n6836;
  assign n6989 = ~n6848 & ~n6988;
  assign n6990 = n6989 ^ n6836;
  assign n6991 = n6837 & ~n6990;
  assign n6992 = n6991 ^ n2583;
  assign n6993 = n6992 ^ n2374;
  assign n6994 = n6633 & ~n6802;
  assign n6995 = n6994 ^ n6635;
  assign n6996 = n6995 ^ n6992;
  assign n6997 = n6993 & n6996;
  assign n6998 = n6997 ^ n2374;
  assign n6999 = n6998 ^ n2194;
  assign n7000 = n6639 & ~n6802;
  assign n7001 = n7000 ^ n6641;
  assign n7002 = n7001 ^ n6998;
  assign n7003 = ~n6999 & ~n7002;
  assign n7004 = n7003 ^ n2194;
  assign n7005 = n6834 & ~n7004;
  assign n7006 = n7005 ^ n6819;
  assign n7007 = n7006 ^ n6819;
  assign n7008 = ~n6831 & ~n7007;
  assign n7009 = n7008 ^ n6819;
  assign n7010 = ~n6820 & ~n7009;
  assign n7011 = n7010 ^ n1621;
  assign n7012 = n7011 ^ n1458;
  assign n7013 = n6662 ^ n1621;
  assign n7014 = ~n6802 & n7013;
  assign n7015 = n7014 ^ n6511;
  assign n7016 = n7015 ^ n7011;
  assign n7017 = n7012 & ~n7016;
  assign n7018 = n7017 ^ n1458;
  assign n7019 = n7018 ^ n1299;
  assign n7020 = n6665 ^ n1458;
  assign n7021 = ~n6802 & n7020;
  assign n7022 = n7021 ^ n6508;
  assign n7023 = n7022 ^ n7018;
  assign n7024 = n7019 & ~n7023;
  assign n7025 = n7024 ^ n1299;
  assign n7026 = n7025 ^ n1158;
  assign n7027 = n6669 & ~n6802;
  assign n7028 = n7027 ^ n6671;
  assign n7029 = n7028 ^ n7025;
  assign n7030 = n7026 & ~n7029;
  assign n7031 = n7030 ^ n1158;
  assign n7032 = n7031 ^ n1027;
  assign n7033 = n6675 & ~n6802;
  assign n7034 = n7033 ^ n6678;
  assign n7035 = n7034 ^ n7031;
  assign n7036 = n7032 & n7035;
  assign n7037 = n7036 ^ n1027;
  assign n7038 = n7037 ^ n905;
  assign n7039 = n6682 & ~n6802;
  assign n7040 = n7039 ^ n6689;
  assign n7041 = n7040 ^ n7037;
  assign n7042 = n7038 & ~n7041;
  assign n7043 = n7042 ^ n905;
  assign n7044 = n7043 ^ n803;
  assign n7045 = n6693 & ~n6802;
  assign n7046 = n7045 ^ n6699;
  assign n7047 = n7046 ^ n7043;
  assign n7048 = n7044 & n7047;
  assign n7049 = n7048 ^ n803;
  assign n7050 = n7049 ^ n707;
  assign n7051 = n6703 & ~n6802;
  assign n7052 = n7051 ^ n6705;
  assign n7053 = n7052 ^ n7049;
  assign n7054 = ~n7050 & ~n7053;
  assign n7055 = n7054 ^ n707;
  assign n7056 = n7055 ^ n608;
  assign n7057 = ~n6709 & ~n6802;
  assign n7058 = n7057 ^ n6711;
  assign n7059 = n7058 ^ n7055;
  assign n7060 = ~n7056 & n7059;
  assign n7061 = n7060 ^ n608;
  assign n7062 = n7061 ^ n514;
  assign n7063 = n6714 ^ n608;
  assign n7064 = ~n6802 & ~n7063;
  assign n7065 = n7064 ^ n6497;
  assign n7066 = n7065 ^ n7061;
  assign n7067 = n7062 & ~n7066;
  assign n7068 = n7067 ^ n514;
  assign n7069 = n7068 ^ n436;
  assign n7070 = n6810 ^ n514;
  assign n7071 = ~n6802 & n7070;
  assign n7072 = n7071 ^ n6494;
  assign n7073 = n7072 ^ n7068;
  assign n7074 = n7069 & n7073;
  assign n7075 = n7074 ^ n436;
  assign n7076 = n7075 ^ n6816;
  assign n7077 = n6817 & ~n7076;
  assign n7078 = n7077 ^ n363;
  assign n7079 = n7078 ^ n6805;
  assign n7080 = ~n6806 & n7079;
  assign n7081 = n7080 ^ n300;
  assign n7082 = n7081 ^ n243;
  assign n7083 = n6729 & ~n6802;
  assign n7084 = n7083 ^ n6735;
  assign n7085 = n7084 ^ n7081;
  assign n7086 = n7082 & ~n7085;
  assign n7087 = n7086 ^ n243;
  assign n7088 = n7087 ^ n210;
  assign n7089 = n6739 & ~n6802;
  assign n7090 = n7089 ^ n6741;
  assign n7091 = n7090 ^ n7087;
  assign n7092 = n7088 & n7091;
  assign n7093 = n7092 ^ n210;
  assign n7094 = n7093 ^ n147;
  assign n7095 = n6745 & ~n6802;
  assign n7096 = n7095 ^ n6748;
  assign n7097 = n7096 ^ n7093;
  assign n7098 = ~n7094 & ~n7097;
  assign n7099 = n7098 ^ n147;
  assign n7100 = n6803 & n7099;
  assign n7101 = n6754 & ~n6760;
  assign n7102 = ~n6802 & ~n7101;
  assign n7103 = n132 & ~n7102;
  assign n7104 = ~n7100 & ~n7103;
  assign n7105 = ~n6486 & ~n7104;
  assign n7106 = ~n6755 & n6757;
  assign n7107 = n7099 & n7106;
  assign n7108 = n132 & n6755;
  assign n7109 = ~n6802 & n7108;
  assign n7110 = ~n7107 & ~n7109;
  assign n7111 = n6760 & ~n6803;
  assign n7112 = ~n7110 & n7111;
  assign n7113 = ~n7105 & ~n7112;
  assign n7114 = n132 & n7099;
  assign n7115 = n6751 ^ n147;
  assign n7116 = ~n6802 & ~n7115;
  assign n7117 = n7116 ^ n6488;
  assign n7118 = ~n7114 & n7117;
  assign n7119 = ~n7113 & ~n7118;
  assign n7120 = n133 & ~n7119;
  assign n7121 = ~n132 & ~n7099;
  assign n7122 = ~n7118 & ~n7121;
  assign n7123 = n6754 ^ n132;
  assign n7124 = ~n6802 & n7123;
  assign n7125 = n7124 ^ n6486;
  assign n7126 = ~n7122 & n7125;
  assign n7127 = n6760 ^ n6758;
  assign n7128 = n6760 ^ n133;
  assign n7129 = n6801 ^ n133;
  assign n7130 = n7129 ^ n133;
  assign n7131 = n7128 & ~n7130;
  assign n7132 = n7131 ^ n133;
  assign n7133 = n7127 & ~n7132;
  assign n7134 = ~n7126 & ~n7133;
  assign n7135 = ~n7120 & n7134;
  assign n7136 = n7078 ^ n300;
  assign n7137 = ~n7135 & n7136;
  assign n7138 = n7137 ^ n6805;
  assign n7139 = n7138 ^ n243;
  assign n7140 = n7075 ^ n363;
  assign n7141 = ~n7135 & n7140;
  assign n7142 = n7141 ^ n6816;
  assign n7143 = n7142 ^ n300;
  assign n7144 = n7019 & ~n7135;
  assign n7145 = n7144 ^ n7022;
  assign n7146 = n7145 ^ n1158;
  assign n7147 = n7012 & ~n7135;
  assign n7148 = n7147 ^ n7015;
  assign n7149 = n7148 ^ n1299;
  assign n7150 = n6993 & ~n7135;
  assign n7151 = n7150 ^ n6995;
  assign n7152 = ~n2194 & ~n7151;
  assign n7153 = ~n6999 & ~n7135;
  assign n7154 = n7153 ^ n7001;
  assign n7155 = n2011 & n7154;
  assign n7156 = ~n7152 & ~n7155;
  assign n7157 = n6954 & ~n7135;
  assign n7158 = n7157 ^ n6956;
  assign n7159 = n7158 ^ n3882;
  assign n7160 = n6950 ^ n4362;
  assign n7161 = ~n7135 & n7160;
  assign n7162 = n7161 ^ n6853;
  assign n7163 = n7162 ^ n4133;
  assign n7164 = n6947 ^ n4606;
  assign n7165 = ~n7135 & n7164;
  assign n7166 = n7165 ^ n6856;
  assign n7167 = n7166 ^ n4362;
  assign n7168 = n6942 & ~n7135;
  assign n7169 = n7168 ^ n6944;
  assign n7170 = n7169 ^ n4606;
  assign n7171 = ~x44 & ~x45;
  assign n7172 = ~x46 & n7171;
  assign n7173 = n6802 & ~n7172;
  assign n7174 = n7135 ^ x47;
  assign n7175 = ~n7173 & n7174;
  assign n7177 = ~n6802 & n7171;
  assign n7176 = ~x47 & ~n7135;
  assign n7178 = n7177 ^ n7176;
  assign n7179 = ~x46 & n7178;
  assign n7180 = n7179 ^ n7176;
  assign n7181 = ~n7175 & ~n7180;
  assign n7182 = n7181 ^ n6479;
  assign n7183 = n6862 ^ n6802;
  assign n7184 = ~n7135 & ~n7183;
  assign n7185 = n7184 ^ n6802;
  assign n7186 = n7185 ^ x48;
  assign n7187 = n7186 ^ n7181;
  assign n7188 = n7182 & n7187;
  assign n7189 = n7188 ^ n6479;
  assign n7190 = n7189 ^ n6181;
  assign n7192 = ~n6864 & n6886;
  assign n7193 = n7192 ^ n6885;
  assign n7194 = n6802 & n7193;
  assign n7195 = n7194 ^ n6885;
  assign n7191 = ~x48 & ~n6802;
  assign n7196 = n7195 ^ n7191;
  assign n7197 = n6862 ^ n6479;
  assign n7198 = n7197 ^ n7195;
  assign n7199 = n7195 ^ n7135;
  assign n7200 = ~n7195 & n7199;
  assign n7201 = n7200 ^ n7195;
  assign n7202 = ~n7198 & ~n7201;
  assign n7203 = n7202 ^ n7200;
  assign n7204 = n7203 ^ n7195;
  assign n7205 = n7204 ^ n7135;
  assign n7206 = n7196 & n7205;
  assign n7207 = n7206 ^ n7191;
  assign n7208 = n7207 ^ x49;
  assign n7209 = n7208 ^ n7189;
  assign n7210 = n7190 & ~n7209;
  assign n7211 = n7210 ^ n6181;
  assign n7212 = n7211 ^ n5905;
  assign n7221 = n6860 ^ x50;
  assign n7213 = n6802 ^ x49;
  assign n7214 = ~n6864 & ~n7213;
  assign n7215 = n6886 & ~n7214;
  assign n7216 = x48 & ~x49;
  assign n7217 = ~n6802 & n7216;
  assign n7218 = ~n7215 & ~n7217;
  assign n7219 = n7218 ^ n6181;
  assign n7220 = ~n7135 & n7219;
  assign n7222 = n7221 ^ n7220;
  assign n7223 = n7222 ^ n7211;
  assign n7224 = n7212 & n7223;
  assign n7225 = n7224 ^ n5905;
  assign n7226 = n7225 ^ n5625;
  assign n7227 = n6920 ^ n5905;
  assign n7228 = n7227 ^ n6901;
  assign n7229 = n7227 & n7228;
  assign n7230 = ~n6899 & n7229;
  assign n7231 = n7230 ^ n7228;
  assign n7232 = n7231 ^ n6920;
  assign n7233 = ~n7135 & ~n7232;
  assign n7234 = n7233 ^ n6920;
  assign n7235 = n7234 ^ n7225;
  assign n7236 = n7226 & ~n7235;
  assign n7237 = n7236 ^ n5625;
  assign n7238 = n7237 ^ n5363;
  assign n7239 = n6924 & ~n7135;
  assign n7240 = n7239 ^ n6926;
  assign n7241 = n7240 ^ n7237;
  assign n7242 = n7238 & n7241;
  assign n7243 = n7242 ^ n5363;
  assign n7244 = n7243 ^ n5108;
  assign n7245 = n6930 & ~n7135;
  assign n7246 = n7245 ^ n6932;
  assign n7247 = n7246 ^ n7243;
  assign n7248 = n7244 & ~n7247;
  assign n7249 = n7248 ^ n5108;
  assign n7250 = n7249 ^ n4851;
  assign n7251 = n6936 & ~n7135;
  assign n7252 = n7251 ^ n6938;
  assign n7253 = n7252 ^ n7249;
  assign n7254 = n7250 & n7253;
  assign n7255 = n7254 ^ n4851;
  assign n7256 = n7255 ^ n7169;
  assign n7257 = n7170 & ~n7256;
  assign n7258 = n7257 ^ n4606;
  assign n7259 = n7258 ^ n7166;
  assign n7260 = ~n7167 & n7259;
  assign n7261 = n7260 ^ n4362;
  assign n7262 = n7261 ^ n7162;
  assign n7263 = n7163 & ~n7262;
  assign n7264 = n7263 ^ n4133;
  assign n7265 = n7264 ^ n7158;
  assign n7266 = ~n7159 & n7265;
  assign n7267 = n7266 ^ n3882;
  assign n7268 = n7267 ^ n3634;
  assign n7269 = n6960 & ~n7135;
  assign n7270 = n7269 ^ n6962;
  assign n7271 = n7270 ^ n7267;
  assign n7272 = ~n7268 & ~n7271;
  assign n7273 = n7272 ^ n3634;
  assign n7274 = n7273 ^ n3397;
  assign n7275 = ~n6966 & ~n7135;
  assign n7276 = n7275 ^ n6969;
  assign n7277 = n7276 ^ n7273;
  assign n7278 = ~n7274 & ~n7277;
  assign n7279 = n7278 ^ n3397;
  assign n7280 = n7279 ^ n3177;
  assign n7281 = ~n6973 & ~n7135;
  assign n7282 = n7281 ^ n6976;
  assign n7283 = n7282 ^ n7279;
  assign n7284 = n7280 & ~n7283;
  assign n7285 = n7284 ^ n3177;
  assign n7286 = n7285 ^ n2980;
  assign n7287 = n6980 & ~n7135;
  assign n7288 = n7287 ^ n6982;
  assign n7289 = n7288 ^ n7285;
  assign n7290 = n7286 & n7289;
  assign n7291 = n7290 ^ n2980;
  assign n7292 = n7291 ^ n2782;
  assign n7293 = n6985 ^ n2980;
  assign n7294 = ~n7135 & n7293;
  assign n7295 = n7294 ^ n6842;
  assign n7296 = n7295 ^ n7291;
  assign n7297 = n7292 & ~n7296;
  assign n7298 = n7297 ^ n2782;
  assign n7299 = n7298 ^ n2583;
  assign n7300 = n6842 ^ n2980;
  assign n7301 = n6985 ^ n6842;
  assign n7302 = n7300 & ~n7301;
  assign n7303 = n7302 ^ n2980;
  assign n7304 = n7303 ^ n2782;
  assign n7305 = ~n7135 & n7304;
  assign n7306 = n7305 ^ n6839;
  assign n7307 = n7306 ^ n7298;
  assign n7308 = n7299 & n7307;
  assign n7309 = n7308 ^ n2583;
  assign n7310 = n7309 ^ n2374;
  assign n7311 = n7303 ^ n6839;
  assign n7312 = ~n6840 & n7311;
  assign n7313 = n7312 ^ n2782;
  assign n7314 = n7313 ^ n2583;
  assign n7315 = ~n7135 & n7314;
  assign n7316 = n7315 ^ n6836;
  assign n7317 = n7316 ^ n7309;
  assign n7318 = n7310 & ~n7317;
  assign n7319 = n7318 ^ n2374;
  assign n7320 = n7156 & ~n7319;
  assign n7321 = n7154 ^ n2011;
  assign n7322 = n2194 & n7151;
  assign n7323 = n7322 ^ n7154;
  assign n7324 = n7321 & n7323;
  assign n7325 = n7324 ^ n2011;
  assign n7326 = ~n7320 & n7325;
  assign n7327 = n7326 ^ n1804;
  assign n7328 = n7004 ^ n2011;
  assign n7329 = ~n7135 & ~n7328;
  assign n7330 = n7329 ^ n6825;
  assign n7331 = n7330 ^ n7326;
  assign n7332 = n7327 & n7331;
  assign n7333 = n7332 ^ n1804;
  assign n7334 = n7333 ^ n1621;
  assign n7335 = n7004 ^ n6825;
  assign n7336 = ~n7328 & ~n7335;
  assign n7337 = n7336 ^ n2011;
  assign n7338 = n7337 ^ n1804;
  assign n7339 = ~n7135 & n7338;
  assign n7340 = n7339 ^ n6822;
  assign n7341 = n7340 ^ n7333;
  assign n7342 = n7334 & ~n7341;
  assign n7343 = n7342 ^ n1621;
  assign n7344 = n7343 ^ n1458;
  assign n7345 = n7337 ^ n6822;
  assign n7346 = n6823 & ~n7345;
  assign n7347 = n7346 ^ n1804;
  assign n7348 = n7347 ^ n1621;
  assign n7349 = ~n7135 & n7348;
  assign n7350 = n7349 ^ n6819;
  assign n7351 = n7350 ^ n7343;
  assign n7352 = n7344 & n7351;
  assign n7353 = n7352 ^ n1458;
  assign n7354 = n7353 ^ n7148;
  assign n7355 = n7149 & ~n7354;
  assign n7356 = n7355 ^ n1299;
  assign n7357 = n7356 ^ n7145;
  assign n7358 = n7146 & ~n7357;
  assign n7359 = n7358 ^ n1158;
  assign n7360 = n7359 ^ n1027;
  assign n7361 = n7026 & ~n7135;
  assign n7362 = n7361 ^ n7028;
  assign n7363 = n7362 ^ n7359;
  assign n7364 = n7360 & ~n7363;
  assign n7365 = n7364 ^ n1027;
  assign n7366 = n7365 ^ n905;
  assign n7367 = n7032 & ~n7135;
  assign n7368 = n7367 ^ n7034;
  assign n7369 = n7368 ^ n7365;
  assign n7370 = n7366 & n7369;
  assign n7371 = n7370 ^ n905;
  assign n7372 = n7371 ^ n803;
  assign n7373 = n7038 & ~n7135;
  assign n7374 = n7373 ^ n7040;
  assign n7375 = n7374 ^ n7371;
  assign n7376 = n7372 & ~n7375;
  assign n7377 = n7376 ^ n803;
  assign n7378 = n7377 ^ n707;
  assign n7379 = n7044 & ~n7135;
  assign n7380 = n7379 ^ n7046;
  assign n7381 = n7380 ^ n7377;
  assign n7382 = ~n7378 & n7381;
  assign n7383 = n7382 ^ n707;
  assign n7384 = n7383 ^ n608;
  assign n7385 = ~n7050 & ~n7135;
  assign n7386 = n7385 ^ n7052;
  assign n7387 = n7386 ^ n7383;
  assign n7388 = ~n7384 & n7387;
  assign n7389 = n7388 ^ n608;
  assign n7390 = n7389 ^ n514;
  assign n7391 = ~n7056 & ~n7135;
  assign n7392 = n7391 ^ n7058;
  assign n7393 = n7392 ^ n7389;
  assign n7394 = n7390 & ~n7393;
  assign n7395 = n7394 ^ n514;
  assign n7396 = n7395 ^ n436;
  assign n7397 = n7062 & ~n7135;
  assign n7398 = n7397 ^ n7065;
  assign n7399 = n7398 ^ n7395;
  assign n7400 = n7396 & ~n7399;
  assign n7401 = n7400 ^ n436;
  assign n7402 = n7401 ^ n363;
  assign n7403 = n7069 & ~n7135;
  assign n7404 = n7403 ^ n7072;
  assign n7405 = n7404 ^ n7401;
  assign n7406 = n7402 & n7405;
  assign n7407 = n7406 ^ n363;
  assign n7408 = n7407 ^ n7142;
  assign n7409 = n7143 & ~n7408;
  assign n7410 = n7409 ^ n300;
  assign n7411 = n7410 ^ n7138;
  assign n7412 = ~n7139 & n7411;
  assign n7413 = n7412 ^ n243;
  assign n7414 = n7413 ^ n210;
  assign n7415 = n7082 & ~n7135;
  assign n7416 = n7415 ^ n7084;
  assign n7417 = n7416 ^ n7413;
  assign n7418 = n7414 & ~n7417;
  assign n7419 = n7418 ^ n210;
  assign n7420 = n7419 ^ n147;
  assign n7421 = n7088 & ~n7135;
  assign n7422 = n7421 ^ n7090;
  assign n7423 = n7422 ^ n7419;
  assign n7424 = ~n7420 & n7423;
  assign n7425 = n7424 ^ n147;
  assign n7426 = n7425 ^ n132;
  assign n7427 = n7099 ^ n132;
  assign n7428 = ~n7135 & n7427;
  assign n7429 = n7428 ^ n7117;
  assign n7430 = ~n133 & ~n7429;
  assign n7431 = ~n7094 & ~n7135;
  assign n7432 = n7431 ^ n7096;
  assign n7433 = n7432 ^ n7425;
  assign n7434 = n7426 & n7433;
  assign n7435 = n7434 ^ n132;
  assign n7436 = ~n7430 & ~n7435;
  assign n7442 = n7118 ^ n7117;
  assign n7443 = ~n7121 & ~n7442;
  assign n7444 = n7443 ^ n7117;
  assign n7445 = ~n7135 & ~n7444;
  assign n7446 = n7445 ^ n7122;
  assign n7447 = n7446 ^ n7445;
  assign n7448 = n7445 ^ n7134;
  assign n7449 = n7448 ^ n7445;
  assign n7450 = ~n7447 & ~n7449;
  assign n7451 = n7450 ^ n7445;
  assign n7452 = ~n133 & ~n7451;
  assign n7453 = n7452 ^ n7445;
  assign n7437 = ~n133 & ~n7122;
  assign n7438 = n1292 & ~n7117;
  assign n7439 = n7099 & n7438;
  assign n7440 = ~n7437 & ~n7439;
  assign n7441 = ~n7135 & ~n7440;
  assign n7454 = n7453 ^ n7441;
  assign n7455 = n7454 ^ n7441;
  assign n7456 = ~n7117 & n7135;
  assign n7457 = n7456 ^ n7441;
  assign n7458 = n7457 ^ n7441;
  assign n7459 = ~n7455 & ~n7458;
  assign n7460 = n7459 ^ n7441;
  assign n7461 = ~n7125 & ~n7460;
  assign n7462 = n7461 ^ n7441;
  assign n7463 = ~n7436 & n7462;
  assign n7464 = n7426 & ~n7463;
  assign n7465 = n7464 ^ n7432;
  assign n7466 = ~n133 & ~n7465;
  assign n7467 = n7407 ^ n300;
  assign n7468 = ~n7463 & n7467;
  assign n7469 = n7468 ^ n7142;
  assign n7470 = n7469 ^ n243;
  assign n7471 = n7402 & ~n7463;
  assign n7472 = n7471 ^ n7404;
  assign n7473 = n7472 ^ n300;
  assign n7474 = n7356 ^ n1158;
  assign n7475 = ~n7463 & n7474;
  assign n7476 = n7475 ^ n7145;
  assign n7477 = n7476 ^ n1027;
  assign n7478 = n7353 ^ n1299;
  assign n7479 = ~n7463 & n7478;
  assign n7480 = n7479 ^ n7148;
  assign n7481 = n7480 ^ n1158;
  assign n7482 = x44 & n7135;
  assign n7483 = ~x42 & ~x43;
  assign n7484 = n7135 & ~n7483;
  assign n7485 = ~n7482 & ~n7484;
  assign n7486 = n7463 ^ x45;
  assign n7487 = n7485 & n7486;
  assign n7489 = ~n7135 & n7483;
  assign n7488 = ~x45 & ~n7463;
  assign n7490 = n7489 ^ n7488;
  assign n7491 = ~x44 & n7490;
  assign n7492 = n7491 ^ n7488;
  assign n7493 = ~n7487 & ~n7492;
  assign n7494 = n7493 ^ n6802;
  assign n7495 = n7171 ^ n7135;
  assign n7496 = ~n7463 & ~n7495;
  assign n7497 = n7496 ^ n7135;
  assign n7498 = n7497 ^ x46;
  assign n7499 = n7498 ^ n7493;
  assign n7500 = n7494 & n7499;
  assign n7501 = n7500 ^ n6802;
  assign n7502 = n7501 ^ n6479;
  assign n7504 = n7172 ^ n6802;
  assign n7505 = n7504 ^ x46;
  assign n7506 = n7505 ^ n7504;
  assign n7507 = n7504 ^ n7172;
  assign n7508 = n7506 & n7507;
  assign n7509 = n7508 ^ n7504;
  assign n7510 = ~n7135 & ~n7509;
  assign n7511 = n7510 ^ n7504;
  assign n7503 = ~x46 & ~n7135;
  assign n7512 = n7511 ^ n7503;
  assign n7513 = n7171 ^ n6802;
  assign n7514 = n7513 ^ n7511;
  assign n7515 = n7511 ^ n7463;
  assign n7516 = n7511 & ~n7515;
  assign n7517 = n7516 ^ n7511;
  assign n7518 = n7514 & n7517;
  assign n7519 = n7518 ^ n7516;
  assign n7520 = n7519 ^ n7511;
  assign n7521 = n7520 ^ n7463;
  assign n7522 = ~n7512 & ~n7521;
  assign n7523 = n7522 ^ n7503;
  assign n7524 = n7523 ^ x47;
  assign n7525 = n7524 ^ n7501;
  assign n7526 = n7502 & ~n7525;
  assign n7527 = n7526 ^ n6479;
  assign n7528 = n7527 ^ n6181;
  assign n7529 = n7182 & ~n7463;
  assign n7530 = n7529 ^ n7186;
  assign n7531 = n7530 ^ n7527;
  assign n7532 = n7528 & n7531;
  assign n7533 = n7532 ^ n6181;
  assign n7534 = n7533 ^ n5905;
  assign n7535 = n7190 & ~n7463;
  assign n7536 = n7535 ^ n7208;
  assign n7537 = n7536 ^ n7533;
  assign n7538 = n7534 & ~n7537;
  assign n7539 = n7538 ^ n5905;
  assign n7540 = n7539 ^ n5625;
  assign n7541 = n7212 & ~n7463;
  assign n7542 = n7541 ^ n7222;
  assign n7543 = n7542 ^ n7539;
  assign n7544 = n7540 & n7543;
  assign n7545 = n7544 ^ n5625;
  assign n7546 = n7545 ^ n5363;
  assign n7547 = n7226 & ~n7463;
  assign n7548 = n7547 ^ n7234;
  assign n7549 = n7548 ^ n7545;
  assign n7550 = n7546 & ~n7549;
  assign n7551 = n7550 ^ n5363;
  assign n7552 = n7551 ^ n5108;
  assign n7553 = n7238 & ~n7463;
  assign n7554 = n7553 ^ n7240;
  assign n7555 = n7554 ^ n7551;
  assign n7556 = n7552 & n7555;
  assign n7557 = n7556 ^ n5108;
  assign n7558 = n7557 ^ n4851;
  assign n7559 = n7244 & ~n7463;
  assign n7560 = n7559 ^ n7246;
  assign n7561 = n7560 ^ n7557;
  assign n7562 = n7558 & ~n7561;
  assign n7563 = n7562 ^ n4851;
  assign n7564 = n7563 ^ n4606;
  assign n7565 = n7250 & ~n7463;
  assign n7566 = n7565 ^ n7252;
  assign n7567 = n7566 ^ n7563;
  assign n7568 = n7564 & n7567;
  assign n7569 = n7568 ^ n4606;
  assign n7570 = n7569 ^ n4362;
  assign n7571 = n7255 ^ n4606;
  assign n7572 = ~n7463 & n7571;
  assign n7573 = n7572 ^ n7169;
  assign n7574 = n7573 ^ n7569;
  assign n7575 = n7570 & ~n7574;
  assign n7576 = n7575 ^ n4362;
  assign n7577 = n7576 ^ n4133;
  assign n7578 = n7258 ^ n4362;
  assign n7579 = ~n7463 & n7578;
  assign n7580 = n7579 ^ n7166;
  assign n7581 = n7580 ^ n7576;
  assign n7582 = n7577 & n7581;
  assign n7583 = n7582 ^ n4133;
  assign n7584 = n7583 ^ n3882;
  assign n7585 = n7261 ^ n4133;
  assign n7586 = ~n7463 & n7585;
  assign n7587 = n7586 ^ n7162;
  assign n7588 = n7587 ^ n7583;
  assign n7589 = n7584 & ~n7588;
  assign n7590 = n7589 ^ n3882;
  assign n7591 = n7590 ^ n3634;
  assign n7592 = n7264 ^ n3882;
  assign n7593 = ~n7463 & n7592;
  assign n7594 = n7593 ^ n7158;
  assign n7595 = n7594 ^ n7590;
  assign n7596 = ~n7591 & n7595;
  assign n7597 = n7596 ^ n3634;
  assign n7598 = n7597 ^ n3397;
  assign n7599 = ~n7268 & ~n7463;
  assign n7600 = n7599 ^ n7270;
  assign n7601 = n7600 ^ n7597;
  assign n7602 = ~n7598 & n7601;
  assign n7603 = n7602 ^ n3397;
  assign n7604 = n7603 ^ n3177;
  assign n7605 = ~n7274 & ~n7463;
  assign n7606 = n7605 ^ n7276;
  assign n7607 = n7606 ^ n7603;
  assign n7608 = n7604 & n7607;
  assign n7609 = n7608 ^ n3177;
  assign n7610 = n7609 ^ n2980;
  assign n7611 = n7280 & ~n7463;
  assign n7612 = n7611 ^ n7282;
  assign n7613 = n7612 ^ n7609;
  assign n7614 = n7610 & ~n7613;
  assign n7615 = n7614 ^ n2980;
  assign n7616 = n7615 ^ n2782;
  assign n7617 = n7286 & ~n7463;
  assign n7618 = n7617 ^ n7288;
  assign n7619 = n7618 ^ n7615;
  assign n7620 = n7616 & n7619;
  assign n7621 = n7620 ^ n2782;
  assign n7622 = n7621 ^ n2583;
  assign n7623 = n7292 & ~n7463;
  assign n7624 = n7623 ^ n7295;
  assign n7625 = n7624 ^ n7621;
  assign n7626 = n7622 & ~n7625;
  assign n7627 = n7626 ^ n2583;
  assign n7628 = n7627 ^ n2374;
  assign n7629 = n7299 & ~n7463;
  assign n7630 = n7629 ^ n7306;
  assign n7631 = n7630 ^ n7627;
  assign n7632 = n7628 & n7631;
  assign n7633 = n7632 ^ n2374;
  assign n7634 = n7633 ^ n2194;
  assign n7635 = n7310 & ~n7463;
  assign n7636 = n7635 ^ n7316;
  assign n7637 = n7636 ^ n7633;
  assign n7638 = ~n7634 & ~n7637;
  assign n7639 = n7638 ^ n2194;
  assign n7640 = n7639 ^ n2011;
  assign n7641 = n7319 ^ n2194;
  assign n7642 = ~n7463 & ~n7641;
  assign n7643 = n7642 ^ n7151;
  assign n7644 = n7643 ^ n7639;
  assign n7645 = ~n7640 & ~n7644;
  assign n7646 = n7645 ^ n2011;
  assign n7647 = n7646 ^ n1804;
  assign n7648 = n7319 ^ n7151;
  assign n7649 = ~n7641 & n7648;
  assign n7650 = n7649 ^ n2194;
  assign n7651 = n7650 ^ n2011;
  assign n7652 = ~n7463 & ~n7651;
  assign n7653 = n7652 ^ n7154;
  assign n7654 = n7653 ^ n7646;
  assign n7655 = n7647 & ~n7654;
  assign n7656 = n7655 ^ n1804;
  assign n7657 = n7656 ^ n1621;
  assign n7658 = n7327 & ~n7463;
  assign n7659 = n7658 ^ n7330;
  assign n7660 = n7659 ^ n7656;
  assign n7661 = n7657 & n7660;
  assign n7662 = n7661 ^ n1621;
  assign n7663 = n7662 ^ n1458;
  assign n7664 = n7334 & ~n7463;
  assign n7665 = n7664 ^ n7340;
  assign n7666 = n7665 ^ n7662;
  assign n7667 = n7663 & ~n7666;
  assign n7668 = n7667 ^ n1458;
  assign n7669 = n7668 ^ n1299;
  assign n7670 = n7344 & ~n7463;
  assign n7671 = n7670 ^ n7350;
  assign n7672 = n7671 ^ n7668;
  assign n7673 = n7669 & n7672;
  assign n7674 = n7673 ^ n1299;
  assign n7675 = n7674 ^ n7480;
  assign n7676 = n7481 & ~n7675;
  assign n7677 = n7676 ^ n1158;
  assign n7678 = n7677 ^ n7476;
  assign n7679 = n7477 & ~n7678;
  assign n7680 = n7679 ^ n1027;
  assign n7681 = n7680 ^ n905;
  assign n7682 = n7360 & ~n7463;
  assign n7683 = n7682 ^ n7362;
  assign n7684 = n7683 ^ n7680;
  assign n7685 = n7681 & ~n7684;
  assign n7686 = n7685 ^ n905;
  assign n7687 = n7686 ^ n803;
  assign n7688 = n7366 & ~n7463;
  assign n7689 = n7688 ^ n7368;
  assign n7690 = n7689 ^ n7686;
  assign n7691 = n7687 & n7690;
  assign n7692 = n7691 ^ n803;
  assign n7693 = n7692 ^ n707;
  assign n7694 = n7372 & ~n7463;
  assign n7695 = n7694 ^ n7374;
  assign n7696 = n7695 ^ n7692;
  assign n7697 = ~n7693 & ~n7696;
  assign n7698 = n7697 ^ n707;
  assign n7699 = n7698 ^ n608;
  assign n7700 = ~n7378 & ~n7463;
  assign n7701 = n7700 ^ n7380;
  assign n7702 = n7701 ^ n7698;
  assign n7703 = ~n7699 & ~n7702;
  assign n7704 = n7703 ^ n608;
  assign n7705 = n7704 ^ n514;
  assign n7706 = ~n7384 & ~n7463;
  assign n7707 = n7706 ^ n7386;
  assign n7708 = n7707 ^ n7704;
  assign n7709 = n7705 & ~n7708;
  assign n7710 = n7709 ^ n514;
  assign n7711 = n7710 ^ n436;
  assign n7712 = n7390 & ~n7463;
  assign n7713 = n7712 ^ n7392;
  assign n7714 = n7713 ^ n7710;
  assign n7715 = n7711 & ~n7714;
  assign n7716 = n7715 ^ n436;
  assign n7717 = n7716 ^ n363;
  assign n7718 = n7396 & ~n7463;
  assign n7719 = n7718 ^ n7398;
  assign n7720 = n7719 ^ n7716;
  assign n7721 = n7717 & ~n7720;
  assign n7722 = n7721 ^ n363;
  assign n7723 = n7722 ^ n7472;
  assign n7724 = ~n7473 & n7723;
  assign n7725 = n7724 ^ n300;
  assign n7726 = n7725 ^ n7469;
  assign n7727 = n7470 & ~n7726;
  assign n7728 = n7727 ^ n243;
  assign n7729 = n7728 ^ n210;
  assign n7730 = n7410 ^ n243;
  assign n7731 = ~n7463 & n7730;
  assign n7732 = n7731 ^ n7138;
  assign n7733 = n7732 ^ n7728;
  assign n7734 = n7729 & n7733;
  assign n7735 = n7734 ^ n210;
  assign n7736 = n7735 ^ n147;
  assign n7737 = n7414 & ~n7463;
  assign n7738 = n7737 ^ n7416;
  assign n7739 = n7738 ^ n7735;
  assign n7740 = ~n7736 & ~n7739;
  assign n7741 = n7740 ^ n147;
  assign n7742 = n7741 ^ n132;
  assign n7743 = ~n7420 & ~n7463;
  assign n7744 = n7743 ^ n7422;
  assign n7745 = n7744 ^ n7741;
  assign n7746 = n7742 & ~n7745;
  assign n7747 = n7746 ^ n132;
  assign n7748 = ~n7466 & ~n7747;
  assign n7749 = ~n7425 & ~n7462;
  assign n7750 = ~n7429 & ~n7462;
  assign n7751 = n133 & ~n7432;
  assign n7752 = ~n7750 & n7751;
  assign n7753 = ~n7749 & n7752;
  assign n7754 = ~n7425 & n7432;
  assign n7755 = n132 & ~n7430;
  assign n7756 = ~n7754 & n7755;
  assign n7757 = ~n7753 & n7756;
  assign n7758 = n7429 ^ n133;
  assign n7759 = n7758 ^ n7429;
  assign n7760 = n129 & ~n7462;
  assign n7761 = n7760 ^ n7429;
  assign n7762 = n7759 & n7761;
  assign n7763 = n7762 ^ n7429;
  assign n7764 = ~n7432 & n7763;
  assign n7765 = n7425 & n7764;
  assign n7766 = ~n7757 & ~n7765;
  assign n7767 = ~n132 & ~n7425;
  assign n7768 = n7767 ^ n7432;
  assign n7769 = n7767 ^ n7429;
  assign n7770 = n7768 & n7769;
  assign n7771 = n7770 ^ n7767;
  assign n7772 = n133 & n7771;
  assign n7773 = n7766 & ~n7772;
  assign n7774 = ~n133 & n7750;
  assign n7775 = ~n7435 & n7774;
  assign n7776 = n7773 & ~n7775;
  assign n7777 = ~n7748 & n7776;
  assign n7778 = x42 & ~n7777;
  assign n7779 = ~x43 & n7778;
  assign n7780 = ~x40 & ~x41;
  assign n7781 = ~x42 & n7780;
  assign n7782 = n7781 ^ n7463;
  assign n7783 = n7777 ^ x43;
  assign n7784 = n7783 ^ n7463;
  assign n7785 = ~n7782 & ~n7784;
  assign n7786 = n7785 ^ n7463;
  assign n7787 = ~n7779 & n7786;
  assign n7788 = n7787 ^ n7135;
  assign n7789 = n7483 ^ n7463;
  assign n7790 = ~n7777 & ~n7789;
  assign n7791 = n7790 ^ n7463;
  assign n7792 = n7791 ^ x44;
  assign n7793 = n7792 ^ n7787;
  assign n7794 = n7788 & n7793;
  assign n7795 = n7794 ^ n7135;
  assign n7796 = n7795 ^ n6802;
  assign n7798 = ~x44 & n7483;
  assign n7799 = n7798 ^ n7135;
  assign n7800 = n7799 ^ n7482;
  assign n7801 = n7463 & ~n7800;
  assign n7802 = n7801 ^ n7482;
  assign n7797 = ~x44 & ~n7463;
  assign n7803 = n7802 ^ n7797;
  assign n7804 = n7483 ^ n7135;
  assign n7805 = n7804 ^ n7802;
  assign n7806 = n7802 ^ n7777;
  assign n7807 = ~n7802 & n7806;
  assign n7808 = n7807 ^ n7802;
  assign n7809 = ~n7805 & ~n7808;
  assign n7810 = n7809 ^ n7807;
  assign n7811 = n7810 ^ n7802;
  assign n7812 = n7811 ^ n7777;
  assign n7813 = n7803 & n7812;
  assign n7814 = n7813 ^ n7797;
  assign n7815 = n7814 ^ x45;
  assign n7816 = n7815 ^ n7795;
  assign n7817 = n7796 & ~n7816;
  assign n7818 = n7817 ^ n6802;
  assign n7819 = n7818 ^ n6479;
  assign n7820 = n7494 & ~n7777;
  assign n7821 = n7820 ^ n7498;
  assign n7822 = n7821 ^ n7818;
  assign n7823 = n7819 & n7822;
  assign n7824 = n7823 ^ n6479;
  assign n7825 = n7824 ^ n6181;
  assign n7826 = n7502 & ~n7777;
  assign n7827 = n7826 ^ n7524;
  assign n7828 = n7827 ^ n7824;
  assign n7829 = n7825 & ~n7828;
  assign n7830 = n7829 ^ n6181;
  assign n7831 = n7830 ^ n5905;
  assign n7832 = n7528 & ~n7777;
  assign n7833 = n7832 ^ n7530;
  assign n7834 = n7833 ^ n7830;
  assign n7835 = n7831 & n7834;
  assign n7836 = n7835 ^ n5905;
  assign n7837 = n7836 ^ n5625;
  assign n7838 = n7534 & ~n7777;
  assign n7839 = n7838 ^ n7536;
  assign n7840 = n7839 ^ n7836;
  assign n7841 = n7837 & ~n7840;
  assign n7842 = n7841 ^ n5625;
  assign n7843 = n7842 ^ n5363;
  assign n7844 = n7540 & ~n7777;
  assign n7845 = n7844 ^ n7542;
  assign n7846 = n7845 ^ n7842;
  assign n7847 = n7843 & n7846;
  assign n7848 = n7847 ^ n5363;
  assign n7849 = n7848 ^ n5108;
  assign n7850 = n7546 & ~n7777;
  assign n7851 = n7850 ^ n7548;
  assign n7852 = n7851 ^ n7848;
  assign n7853 = n7849 & ~n7852;
  assign n7854 = n7853 ^ n5108;
  assign n7855 = n7854 ^ n4851;
  assign n7856 = n7552 & ~n7777;
  assign n7857 = n7856 ^ n7554;
  assign n7858 = n7857 ^ n7854;
  assign n7859 = n7855 & n7858;
  assign n7860 = n7859 ^ n4851;
  assign n7861 = n7860 ^ n4606;
  assign n7862 = n7742 & ~n7777;
  assign n7863 = n7862 ^ n7744;
  assign n7864 = ~n133 & n7863;
  assign n7865 = n7705 & ~n7777;
  assign n7866 = n7865 ^ n7707;
  assign n7867 = n7866 ^ n436;
  assign n7868 = ~n7699 & ~n7777;
  assign n7869 = n7868 ^ n7701;
  assign n7870 = n7869 ^ n514;
  assign n7871 = n7584 & ~n7777;
  assign n7872 = n7871 ^ n7587;
  assign n7873 = n7872 ^ n3634;
  assign n7874 = n7577 & ~n7777;
  assign n7875 = n7874 ^ n7580;
  assign n7876 = n7875 ^ n3882;
  assign n7877 = n7558 & ~n7777;
  assign n7878 = n7877 ^ n7560;
  assign n7879 = n7878 ^ n7860;
  assign n7880 = n7861 & ~n7879;
  assign n7881 = n7880 ^ n4606;
  assign n7882 = n7881 ^ n4362;
  assign n7883 = n7564 & ~n7777;
  assign n7884 = n7883 ^ n7566;
  assign n7885 = n7884 ^ n7881;
  assign n7886 = n7882 & n7885;
  assign n7887 = n7886 ^ n4362;
  assign n7888 = n7887 ^ n4133;
  assign n7889 = n7570 & ~n7777;
  assign n7890 = n7889 ^ n7573;
  assign n7891 = n7890 ^ n7887;
  assign n7892 = n7888 & ~n7891;
  assign n7893 = n7892 ^ n4133;
  assign n7894 = n7893 ^ n7875;
  assign n7895 = ~n7876 & n7894;
  assign n7896 = n7895 ^ n3882;
  assign n7897 = n7896 ^ n7872;
  assign n7898 = ~n7873 & ~n7897;
  assign n7899 = n7898 ^ n3634;
  assign n7900 = n7899 ^ n3397;
  assign n7901 = ~n7591 & ~n7777;
  assign n7902 = n7901 ^ n7594;
  assign n7903 = n7902 ^ n7899;
  assign n7904 = ~n7900 & ~n7903;
  assign n7905 = n7904 ^ n3397;
  assign n7906 = n7905 ^ n3177;
  assign n7907 = ~n7598 & ~n7777;
  assign n7908 = n7907 ^ n7600;
  assign n7909 = n7908 ^ n7905;
  assign n7910 = n7906 & ~n7909;
  assign n7911 = n7910 ^ n3177;
  assign n7912 = n7911 ^ n2980;
  assign n7913 = n7604 & ~n7777;
  assign n7914 = n7913 ^ n7606;
  assign n7915 = n7914 ^ n7911;
  assign n7916 = n7912 & n7915;
  assign n7917 = n7916 ^ n2980;
  assign n7918 = n7917 ^ n2782;
  assign n7919 = n7610 & ~n7777;
  assign n7920 = n7919 ^ n7612;
  assign n7921 = n7920 ^ n7917;
  assign n7922 = n7918 & ~n7921;
  assign n7923 = n7922 ^ n2782;
  assign n7924 = n7923 ^ n2583;
  assign n7925 = n7616 & ~n7777;
  assign n7926 = n7925 ^ n7618;
  assign n7927 = n7926 ^ n7923;
  assign n7928 = n7924 & n7927;
  assign n7929 = n7928 ^ n2583;
  assign n7930 = n7929 ^ n2374;
  assign n7931 = n7622 & ~n7777;
  assign n7932 = n7931 ^ n7624;
  assign n7933 = n7932 ^ n7929;
  assign n7934 = n7930 & ~n7933;
  assign n7935 = n7934 ^ n2374;
  assign n7936 = n7935 ^ n2194;
  assign n7937 = n7628 & ~n7777;
  assign n7938 = n7937 ^ n7630;
  assign n7939 = n7938 ^ n7935;
  assign n7940 = ~n7936 & n7939;
  assign n7941 = n7940 ^ n2194;
  assign n7942 = n7941 ^ n2011;
  assign n7943 = ~n7634 & ~n7777;
  assign n7944 = n7943 ^ n7636;
  assign n7945 = n7944 ^ n7941;
  assign n7946 = ~n7942 & n7945;
  assign n7947 = n7946 ^ n2011;
  assign n7948 = n7947 ^ n1804;
  assign n7949 = ~n7640 & ~n7777;
  assign n7950 = n7949 ^ n7643;
  assign n7951 = n7950 ^ n7947;
  assign n7952 = n7948 & n7951;
  assign n7953 = n7952 ^ n1804;
  assign n7954 = n7953 ^ n1621;
  assign n7955 = n7647 & ~n7777;
  assign n7956 = n7955 ^ n7653;
  assign n7957 = n7956 ^ n7953;
  assign n7958 = n7954 & ~n7957;
  assign n7959 = n7958 ^ n1621;
  assign n7960 = n7959 ^ n1458;
  assign n7961 = n7657 & ~n7777;
  assign n7962 = n7961 ^ n7659;
  assign n7963 = n7962 ^ n7959;
  assign n7964 = n7960 & n7963;
  assign n7965 = n7964 ^ n1458;
  assign n7966 = n7965 ^ n1299;
  assign n7967 = n7663 & ~n7777;
  assign n7968 = n7967 ^ n7665;
  assign n7969 = n7968 ^ n7965;
  assign n7970 = n7966 & ~n7969;
  assign n7971 = n7970 ^ n1299;
  assign n7972 = n7971 ^ n1158;
  assign n7973 = n7669 & ~n7777;
  assign n7974 = n7973 ^ n7671;
  assign n7975 = n7974 ^ n7971;
  assign n7976 = n7972 & n7975;
  assign n7977 = n7976 ^ n1158;
  assign n7978 = n7977 ^ n1027;
  assign n7979 = n7674 ^ n1158;
  assign n7980 = ~n7777 & n7979;
  assign n7981 = n7980 ^ n7480;
  assign n7982 = n7981 ^ n7977;
  assign n7983 = n7978 & ~n7982;
  assign n7984 = n7983 ^ n1027;
  assign n7985 = n7984 ^ n905;
  assign n7986 = n7677 ^ n1027;
  assign n7987 = ~n7777 & n7986;
  assign n7988 = n7987 ^ n7476;
  assign n7989 = n7988 ^ n7984;
  assign n7990 = n7985 & ~n7989;
  assign n7991 = n7990 ^ n905;
  assign n7992 = n7991 ^ n803;
  assign n7993 = n7681 & ~n7777;
  assign n7994 = n7993 ^ n7683;
  assign n7995 = n7994 ^ n7991;
  assign n7996 = n7992 & ~n7995;
  assign n7997 = n7996 ^ n803;
  assign n7998 = n7997 ^ n707;
  assign n7999 = n7687 & ~n7777;
  assign n8000 = n7999 ^ n7689;
  assign n8001 = n8000 ^ n7997;
  assign n8002 = ~n7998 & n8001;
  assign n8003 = n8002 ^ n707;
  assign n8004 = n8003 ^ n608;
  assign n8005 = ~n7693 & ~n7777;
  assign n8006 = n8005 ^ n7695;
  assign n8007 = n8006 ^ n8003;
  assign n8008 = ~n8004 & n8007;
  assign n8009 = n8008 ^ n608;
  assign n8010 = n8009 ^ n7869;
  assign n8011 = ~n7870 & n8010;
  assign n8012 = n8011 ^ n514;
  assign n8013 = n8012 ^ n7866;
  assign n8014 = n7867 & ~n8013;
  assign n8015 = n8014 ^ n436;
  assign n8016 = n8015 ^ n363;
  assign n8017 = n7711 & ~n7777;
  assign n8018 = n8017 ^ n7713;
  assign n8019 = n8018 ^ n8015;
  assign n8020 = n8016 & ~n8019;
  assign n8021 = n8020 ^ n363;
  assign n8022 = n8021 ^ n300;
  assign n8023 = n7717 & ~n7777;
  assign n8024 = n8023 ^ n7719;
  assign n8025 = n8024 ^ n8021;
  assign n8026 = n8022 & ~n8025;
  assign n8027 = n8026 ^ n300;
  assign n8028 = n8027 ^ n243;
  assign n8029 = n7722 ^ n300;
  assign n8030 = ~n7777 & n8029;
  assign n8031 = n8030 ^ n7472;
  assign n8032 = n8031 ^ n8027;
  assign n8033 = n8028 & n8032;
  assign n8034 = n8033 ^ n243;
  assign n8035 = n8034 ^ n210;
  assign n8036 = n7725 ^ n243;
  assign n8037 = ~n7777 & n8036;
  assign n8038 = n8037 ^ n7469;
  assign n8039 = n8038 ^ n8034;
  assign n8040 = n8035 & ~n8039;
  assign n8041 = n8040 ^ n210;
  assign n8042 = n8041 ^ n147;
  assign n8043 = n7729 & ~n7777;
  assign n8044 = n8043 ^ n7732;
  assign n8045 = n8044 ^ n8041;
  assign n8046 = ~n8042 & n8045;
  assign n8047 = n8046 ^ n147;
  assign n8048 = n8047 ^ n132;
  assign n8049 = ~n7736 & ~n7777;
  assign n8050 = n8049 ^ n7738;
  assign n8051 = n8050 ^ n8047;
  assign n8052 = n8048 & n8051;
  assign n8053 = n8052 ^ n132;
  assign n8054 = ~n7864 & ~n8053;
  assign n8055 = ~n7465 & ~n7776;
  assign n8056 = ~n7747 & n8055;
  assign n8057 = ~n7741 & ~n7744;
  assign n8058 = n132 & n7465;
  assign n8059 = ~n8057 & n8058;
  assign n8060 = ~n133 & ~n8059;
  assign n8061 = ~n8056 & n8060;
  assign n8062 = n7744 & ~n7776;
  assign n8063 = n7741 & n8062;
  assign n8064 = ~n7465 & ~n8063;
  assign n8065 = n132 & ~n7776;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~n132 & ~n7744;
  assign n8068 = ~n7465 & ~n8067;
  assign n8069 = ~n7741 & ~n8068;
  assign n8070 = n133 & ~n8069;
  assign n8071 = n7745 ^ n7741;
  assign n8072 = n8055 ^ n7741;
  assign n8073 = n8071 & n8072;
  assign n8074 = n8073 ^ n7741;
  assign n8075 = n132 & n8074;
  assign n8076 = n8070 & ~n8075;
  assign n8077 = ~n8066 & n8076;
  assign n8078 = ~n8061 & ~n8077;
  assign n8079 = ~n132 & n7741;
  assign n8080 = n7465 & n7744;
  assign n8081 = n8079 & n8080;
  assign n8082 = ~n8078 & ~n8081;
  assign n8083 = ~n8054 & n8082;
  assign n8084 = n7861 & ~n8083;
  assign n8085 = n8084 ^ n7878;
  assign n8086 = ~n4362 & ~n8085;
  assign n8087 = n7882 & ~n8083;
  assign n8088 = n8087 ^ n7884;
  assign n8089 = ~n4133 & n8088;
  assign n8090 = ~n8086 & ~n8089;
  assign n8091 = n7788 & ~n8083;
  assign n8092 = n8091 ^ n7792;
  assign n8093 = n8092 ^ n6802;
  assign n8094 = ~x38 & ~x39;
  assign n8095 = ~x40 & n8094;
  assign n8096 = x41 & ~n8095;
  assign n8097 = ~n8083 & ~n8096;
  assign n8098 = n7780 & n8094;
  assign n8099 = x42 & ~n8098;
  assign n8100 = n7777 & n8099;
  assign n8101 = ~n8097 & n8100;
  assign n8102 = ~n7777 & n8095;
  assign n8103 = n7780 & ~n8102;
  assign n8104 = n8103 ^ n8083;
  assign n8105 = n8104 ^ n8103;
  assign n8106 = ~n7777 & n8096;
  assign n8107 = n8106 ^ n8103;
  assign n8108 = n8105 & n8107;
  assign n8109 = n8108 ^ n8103;
  assign n8110 = ~x42 & n8109;
  assign n8111 = ~n8101 & ~n8110;
  assign n8112 = ~n7463 & n8111;
  assign n8113 = ~n7780 & ~n8083;
  assign n8114 = n7777 & ~n8095;
  assign n8115 = x41 & n8114;
  assign n8116 = n8113 & ~n8115;
  assign n8117 = n7777 & n8083;
  assign n8118 = n8098 & n8117;
  assign n8119 = ~n8116 & ~n8118;
  assign n8120 = ~x42 & ~n8119;
  assign n8121 = ~n8083 & ~n8098;
  assign n8122 = n7778 & ~n8096;
  assign n8123 = ~n8121 & n8122;
  assign n8124 = ~n8120 & ~n8123;
  assign n8125 = ~n8112 & n8124;
  assign n8126 = n8125 ^ n7135;
  assign n8128 = n7777 ^ n7463;
  assign n8129 = n8128 ^ n7777;
  assign n8130 = n8129 ^ n8128;
  assign n8131 = n8128 ^ n7780;
  assign n8132 = n8130 & n8131;
  assign n8133 = n8132 ^ n8128;
  assign n8134 = ~x42 & n8133;
  assign n8135 = n8134 ^ n8128;
  assign n8127 = ~x42 & ~n7777;
  assign n8136 = n8135 ^ n8127;
  assign n8137 = n7780 ^ n7463;
  assign n8138 = n8137 ^ n8135;
  assign n8139 = n8135 ^ n8083;
  assign n8140 = ~n8135 & n8139;
  assign n8141 = n8140 ^ n8135;
  assign n8142 = ~n8138 & ~n8141;
  assign n8143 = n8142 ^ n8140;
  assign n8144 = n8143 ^ n8135;
  assign n8145 = n8144 ^ n8083;
  assign n8146 = n8136 & n8145;
  assign n8147 = n8146 ^ n8127;
  assign n8148 = n8147 ^ x43;
  assign n8149 = n8148 ^ n8125;
  assign n8150 = n8126 & ~n8149;
  assign n8151 = n8150 ^ n7135;
  assign n8152 = n8151 ^ n8092;
  assign n8153 = ~n8093 & n8152;
  assign n8154 = n8153 ^ n6802;
  assign n8155 = n8154 ^ n6479;
  assign n8156 = n7796 & ~n8083;
  assign n8157 = n8156 ^ n7815;
  assign n8158 = n8157 ^ n8154;
  assign n8159 = n8155 & ~n8158;
  assign n8160 = n8159 ^ n6479;
  assign n8161 = n8160 ^ n6181;
  assign n8162 = n7819 & ~n8083;
  assign n8163 = n8162 ^ n7821;
  assign n8164 = n8163 ^ n8160;
  assign n8165 = n8161 & n8164;
  assign n8166 = n8165 ^ n6181;
  assign n8167 = n8166 ^ n5905;
  assign n8168 = n7825 & ~n8083;
  assign n8169 = n8168 ^ n7827;
  assign n8170 = n8169 ^ n8166;
  assign n8171 = n8167 & ~n8170;
  assign n8172 = n8171 ^ n5905;
  assign n8173 = n8172 ^ n5625;
  assign n8174 = n7831 & ~n8083;
  assign n8175 = n8174 ^ n7833;
  assign n8176 = n8175 ^ n8172;
  assign n8177 = n8173 & n8176;
  assign n8178 = n8177 ^ n5625;
  assign n8179 = n8178 ^ n5363;
  assign n8180 = n7837 & ~n8083;
  assign n8181 = n8180 ^ n7839;
  assign n8182 = n8181 ^ n8178;
  assign n8183 = n8179 & ~n8182;
  assign n8184 = n8183 ^ n5363;
  assign n8185 = n8184 ^ n5108;
  assign n8186 = n7843 & ~n8083;
  assign n8187 = n8186 ^ n7845;
  assign n8188 = n8187 ^ n8184;
  assign n8189 = n8185 & n8188;
  assign n8190 = n8189 ^ n5108;
  assign n8191 = n8190 ^ n4851;
  assign n8192 = n7849 & ~n8083;
  assign n8193 = n8192 ^ n7851;
  assign n8194 = n8193 ^ n8190;
  assign n8195 = n8191 & ~n8194;
  assign n8196 = n8195 ^ n4851;
  assign n8197 = n8196 ^ n4606;
  assign n8198 = n7855 & ~n8083;
  assign n8199 = n8198 ^ n7857;
  assign n8200 = n8199 ^ n8196;
  assign n8201 = n8197 & n8200;
  assign n8202 = n8201 ^ n4606;
  assign n8203 = n8090 & n8202;
  assign n8204 = n8088 ^ n4133;
  assign n8205 = n4362 & n8085;
  assign n8206 = n8205 ^ n8088;
  assign n8207 = ~n8204 & n8206;
  assign n8208 = n8207 ^ n4133;
  assign n8209 = ~n8203 & ~n8208;
  assign n8210 = n8209 ^ n3882;
  assign n8211 = n7888 & ~n8083;
  assign n8212 = n8211 ^ n7890;
  assign n8213 = n8212 ^ n8209;
  assign n8214 = ~n8210 & n8213;
  assign n8215 = n8214 ^ n3882;
  assign n8216 = n8215 ^ n3634;
  assign n8217 = n7893 ^ n3882;
  assign n8218 = ~n8083 & n8217;
  assign n8219 = n8218 ^ n7875;
  assign n8220 = n8219 ^ n8215;
  assign n8221 = ~n8216 & n8220;
  assign n8222 = n8221 ^ n3634;
  assign n8223 = n8222 ^ n3397;
  assign n8224 = n7896 ^ n3634;
  assign n8225 = ~n8083 & ~n8224;
  assign n8226 = n8225 ^ n7872;
  assign n8227 = n8226 ^ n8222;
  assign n8228 = ~n8223 & n8227;
  assign n8229 = n8228 ^ n3397;
  assign n8230 = n8229 ^ n3177;
  assign n8231 = ~n7900 & ~n8083;
  assign n8232 = n8231 ^ n7902;
  assign n8233 = n8232 ^ n8229;
  assign n8234 = n8230 & n8233;
  assign n8235 = n8234 ^ n3177;
  assign n8236 = n8235 ^ n2980;
  assign n8237 = n7906 & ~n8083;
  assign n8238 = n8237 ^ n7908;
  assign n8239 = n8238 ^ n8235;
  assign n8240 = n8236 & ~n8239;
  assign n8241 = n8240 ^ n2980;
  assign n8242 = n8241 ^ n2782;
  assign n8243 = n7912 & ~n8083;
  assign n8244 = n8243 ^ n7914;
  assign n8245 = n8244 ^ n8241;
  assign n8246 = n8242 & n8245;
  assign n8247 = n8246 ^ n2782;
  assign n8248 = n8247 ^ n2583;
  assign n8249 = n7918 & ~n8083;
  assign n8250 = n8249 ^ n7920;
  assign n8251 = n8250 ^ n8247;
  assign n8252 = n8248 & ~n8251;
  assign n8253 = n8252 ^ n2583;
  assign n8254 = n8253 ^ n2374;
  assign n8255 = n8048 & ~n8083;
  assign n8256 = n8255 ^ n8050;
  assign n8257 = ~n133 & ~n8256;
  assign n8258 = n8022 & ~n8083;
  assign n8259 = n8258 ^ n8024;
  assign n8260 = n8259 ^ n243;
  assign n8261 = n8016 & ~n8083;
  assign n8262 = n8261 ^ n8018;
  assign n8263 = n8262 ^ n300;
  assign n8264 = n8012 ^ n436;
  assign n8265 = ~n8083 & n8264;
  assign n8266 = n8265 ^ n7866;
  assign n8267 = n8266 ^ n363;
  assign n8268 = ~n7998 & ~n8083;
  assign n8269 = n8268 ^ n8000;
  assign n8270 = n8269 ^ n608;
  assign n8271 = n7992 & ~n8083;
  assign n8272 = n8271 ^ n7994;
  assign n8273 = n8272 ^ n707;
  assign n8274 = n7985 & ~n8083;
  assign n8275 = n8274 ^ n7988;
  assign n8276 = n803 & n8275;
  assign n8277 = n8276 ^ n8272;
  assign n8278 = ~n8273 & n8277;
  assign n8279 = n8278 ^ n8272;
  assign n8280 = n8279 ^ n8269;
  assign n8281 = n8280 ^ n8269;
  assign n8282 = ~n803 & ~n8275;
  assign n8283 = n707 & ~n8272;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = n7924 & ~n8083;
  assign n8286 = n8285 ^ n7926;
  assign n8287 = n8286 ^ n8253;
  assign n8288 = n8254 & n8287;
  assign n8289 = n8288 ^ n2374;
  assign n8290 = n8289 ^ n2194;
  assign n8291 = n7930 & ~n8083;
  assign n8292 = n8291 ^ n7932;
  assign n8293 = n8292 ^ n8289;
  assign n8294 = ~n8290 & ~n8293;
  assign n8295 = n8294 ^ n2194;
  assign n8296 = n8295 ^ n2011;
  assign n8297 = ~n7936 & ~n8083;
  assign n8298 = n8297 ^ n7938;
  assign n8299 = n8298 ^ n8295;
  assign n8300 = ~n8296 & ~n8299;
  assign n8301 = n8300 ^ n2011;
  assign n8302 = n8301 ^ n1804;
  assign n8303 = ~n7942 & ~n8083;
  assign n8304 = n8303 ^ n7944;
  assign n8305 = n8304 ^ n8301;
  assign n8306 = n8302 & ~n8305;
  assign n8307 = n8306 ^ n1804;
  assign n8308 = n8307 ^ n1621;
  assign n8309 = n7948 & ~n8083;
  assign n8310 = n8309 ^ n7950;
  assign n8311 = n8310 ^ n8307;
  assign n8312 = n8308 & n8311;
  assign n8313 = n8312 ^ n1621;
  assign n8314 = n8313 ^ n1458;
  assign n8315 = n7954 & ~n8083;
  assign n8316 = n8315 ^ n7956;
  assign n8317 = n8316 ^ n8313;
  assign n8318 = n8314 & ~n8317;
  assign n8319 = n8318 ^ n1458;
  assign n8320 = n8319 ^ n1299;
  assign n8321 = n7960 & ~n8083;
  assign n8322 = n8321 ^ n7962;
  assign n8323 = n8322 ^ n8319;
  assign n8324 = n8320 & n8323;
  assign n8325 = n8324 ^ n1299;
  assign n8326 = n8325 ^ n1158;
  assign n8327 = n7966 & ~n8083;
  assign n8328 = n8327 ^ n7968;
  assign n8329 = n8328 ^ n8325;
  assign n8330 = n8326 & ~n8329;
  assign n8331 = n8330 ^ n1158;
  assign n8332 = n8331 ^ n1027;
  assign n8333 = n7972 & ~n8083;
  assign n8334 = n8333 ^ n7974;
  assign n8335 = n8334 ^ n8331;
  assign n8336 = n8332 & n8335;
  assign n8337 = n8336 ^ n1027;
  assign n8338 = n8337 ^ n905;
  assign n8339 = n7978 & ~n8083;
  assign n8340 = n8339 ^ n7981;
  assign n8341 = n8340 ^ n8337;
  assign n8342 = n8338 & ~n8341;
  assign n8343 = n8342 ^ n905;
  assign n8344 = n8284 & n8343;
  assign n8345 = n8344 ^ n8269;
  assign n8346 = n8345 ^ n8269;
  assign n8347 = ~n8281 & ~n8346;
  assign n8348 = n8347 ^ n8269;
  assign n8349 = ~n8270 & ~n8348;
  assign n8350 = n8349 ^ n608;
  assign n8351 = n8350 ^ n514;
  assign n8352 = ~n8004 & ~n8083;
  assign n8353 = n8352 ^ n8006;
  assign n8354 = n8353 ^ n8350;
  assign n8355 = n8351 & ~n8354;
  assign n8356 = n8355 ^ n514;
  assign n8357 = n8356 ^ n436;
  assign n8358 = n8009 ^ n514;
  assign n8359 = ~n8083 & n8358;
  assign n8360 = n8359 ^ n7869;
  assign n8361 = n8360 ^ n8356;
  assign n8362 = n8357 & n8361;
  assign n8363 = n8362 ^ n436;
  assign n8364 = n8363 ^ n8266;
  assign n8365 = n8267 & ~n8364;
  assign n8366 = n8365 ^ n363;
  assign n8367 = n8366 ^ n8262;
  assign n8368 = n8263 & ~n8367;
  assign n8369 = n8368 ^ n300;
  assign n8370 = n8369 ^ n8259;
  assign n8371 = n8260 & ~n8370;
  assign n8372 = n8371 ^ n243;
  assign n8373 = n8372 ^ n210;
  assign n8374 = n8028 & ~n8083;
  assign n8375 = n8374 ^ n8031;
  assign n8376 = n8375 ^ n8372;
  assign n8377 = n8373 & n8376;
  assign n8378 = n8377 ^ n210;
  assign n8379 = n8378 ^ n147;
  assign n8380 = n8035 & ~n8083;
  assign n8381 = n8380 ^ n8038;
  assign n8382 = n8381 ^ n8378;
  assign n8383 = ~n8379 & ~n8382;
  assign n8384 = n8383 ^ n147;
  assign n8385 = n8384 ^ n132;
  assign n8386 = ~n8042 & ~n8083;
  assign n8387 = n8386 ^ n8044;
  assign n8388 = n8387 ^ n8384;
  assign n8389 = n8385 & ~n8388;
  assign n8390 = n8389 ^ n132;
  assign n8391 = ~n8257 & ~n8390;
  assign n8392 = n7863 & n8053;
  assign n8393 = n7863 & ~n8082;
  assign n8394 = n8050 & ~n8393;
  assign n8395 = n8394 ^ n8047;
  assign n8396 = n8394 ^ n7863;
  assign n8397 = n8394 ^ n8048;
  assign n8398 = ~n8394 & n8397;
  assign n8399 = n8398 ^ n8394;
  assign n8400 = ~n8396 & ~n8399;
  assign n8401 = n8400 ^ n8398;
  assign n8402 = n8401 ^ n8394;
  assign n8403 = n8402 ^ n8048;
  assign n8404 = ~n8395 & n8403;
  assign n8405 = n8404 ^ n8394;
  assign n8406 = ~n8392 & ~n8405;
  assign n8407 = ~n133 & ~n8406;
  assign n8408 = n7863 & n8082;
  assign n8409 = ~n8050 & n8408;
  assign n8410 = ~n132 & n8051;
  assign n8411 = n133 & ~n8410;
  assign n8412 = n8047 & ~n8050;
  assign n8413 = ~n8082 & n8412;
  assign n8414 = n8413 ^ n7863;
  assign n8415 = n8414 ^ n8413;
  assign n8416 = n8413 ^ n8053;
  assign n8417 = n8415 & ~n8416;
  assign n8418 = n8417 ^ n8413;
  assign n8419 = n8411 & n8418;
  assign n8420 = ~n8409 & ~n8419;
  assign n8421 = ~n8407 & n8420;
  assign n8422 = ~n8391 & ~n8421;
  assign n8423 = n8254 & ~n8422;
  assign n8424 = n8423 ^ n8286;
  assign n8425 = n8424 ^ n2194;
  assign n8426 = n8248 & ~n8422;
  assign n8427 = n8426 ^ n8250;
  assign n8428 = n8427 ^ n2374;
  assign n8429 = n8236 & ~n8422;
  assign n8430 = n8429 ^ n8238;
  assign n8431 = n8430 ^ n2782;
  assign n8432 = n8230 & ~n8422;
  assign n8433 = n8432 ^ n8232;
  assign n8434 = n8433 ^ n2980;
  assign n8435 = n8179 & ~n8422;
  assign n8436 = n8435 ^ n8181;
  assign n8437 = n8436 ^ n5108;
  assign n8438 = n8173 & ~n8422;
  assign n8439 = n8438 ^ n8175;
  assign n8440 = n8439 ^ n5363;
  assign n8441 = n8151 ^ n6802;
  assign n8442 = ~n8422 & n8441;
  assign n8443 = n8442 ^ n8092;
  assign n8444 = n8443 ^ n6479;
  assign n8457 = ~n8113 & ~n8117;
  assign n8458 = n8457 ^ x42;
  assign n8445 = n8095 ^ n7777;
  assign n8446 = n8095 ^ x41;
  assign n8447 = n8446 ^ n8095;
  assign n8448 = n8095 ^ n8083;
  assign n8449 = n8448 ^ n8095;
  assign n8450 = ~n8447 & n8449;
  assign n8451 = n8450 ^ n8095;
  assign n8452 = ~n8445 & ~n8451;
  assign n8453 = n8452 ^ n7777;
  assign n8454 = ~n8116 & n8453;
  assign n8455 = n8454 ^ n7463;
  assign n8456 = ~n8422 & n8455;
  assign n8459 = n8458 ^ n8456;
  assign n8460 = n7135 & n8459;
  assign n8461 = x38 & ~n8422;
  assign n8462 = ~x39 & n8461;
  assign n8463 = ~x36 & ~x37;
  assign n8464 = ~x38 & n8463;
  assign n8465 = n8464 ^ n8083;
  assign n8466 = n8422 ^ x39;
  assign n8467 = n8466 ^ n8083;
  assign n8468 = ~n8465 & ~n8467;
  assign n8469 = n8468 ^ n8083;
  assign n8470 = ~n8462 & n8469;
  assign n8471 = n8470 ^ n7777;
  assign n8472 = n8094 ^ n8083;
  assign n8473 = ~n8422 & ~n8472;
  assign n8474 = n8473 ^ n8083;
  assign n8475 = n8474 ^ x40;
  assign n8476 = n8475 ^ n8470;
  assign n8477 = n8471 & n8476;
  assign n8478 = n8477 ^ n7777;
  assign n8479 = n8478 ^ n7463;
  assign n8481 = x40 & n7777;
  assign n8482 = n8481 ^ n8445;
  assign n8483 = ~n8083 & ~n8482;
  assign n8484 = n8483 ^ n8445;
  assign n8480 = ~x40 & ~n8083;
  assign n8485 = n8484 ^ n8480;
  assign n8486 = n8094 ^ n7777;
  assign n8487 = n8486 ^ n8484;
  assign n8488 = n8484 ^ n8422;
  assign n8489 = n8484 & ~n8488;
  assign n8490 = n8489 ^ n8484;
  assign n8491 = n8487 & n8490;
  assign n8492 = n8491 ^ n8489;
  assign n8493 = n8492 ^ n8484;
  assign n8494 = n8493 ^ n8422;
  assign n8495 = ~n8485 & ~n8494;
  assign n8496 = n8495 ^ n8480;
  assign n8497 = n8496 ^ x41;
  assign n8498 = n8497 ^ n8478;
  assign n8499 = n8479 & ~n8498;
  assign n8500 = n8499 ^ n7463;
  assign n8501 = ~n8460 & ~n8500;
  assign n8502 = ~n7135 & ~n8459;
  assign n8503 = ~n8111 & ~n8125;
  assign n8504 = ~n8126 & n8503;
  assign n8505 = n8504 ^ n8126;
  assign n8506 = ~n8422 & n8505;
  assign n8507 = n8506 ^ n8148;
  assign n8508 = ~n8502 & n8507;
  assign n8509 = ~n8501 & n8508;
  assign n8510 = ~n6802 & ~n8509;
  assign n8511 = n8510 ^ n8443;
  assign n8512 = n8511 ^ n8443;
  assign n8513 = ~n8501 & ~n8502;
  assign n8514 = ~n8507 & ~n8513;
  assign n8515 = n8514 ^ n8443;
  assign n8516 = n8515 ^ n8443;
  assign n8517 = ~n8512 & ~n8516;
  assign n8518 = n8517 ^ n8443;
  assign n8519 = ~n8444 & n8518;
  assign n8520 = n8519 ^ n6479;
  assign n8521 = n8520 ^ n6181;
  assign n8522 = n8155 & ~n8422;
  assign n8523 = n8522 ^ n8157;
  assign n8524 = n8523 ^ n8520;
  assign n8525 = n8521 & ~n8524;
  assign n8526 = n8525 ^ n6181;
  assign n8527 = n8526 ^ n5905;
  assign n8528 = n8161 & ~n8422;
  assign n8529 = n8528 ^ n8163;
  assign n8530 = n8529 ^ n8526;
  assign n8531 = n8527 & n8530;
  assign n8532 = n8531 ^ n5905;
  assign n8533 = n8532 ^ n5625;
  assign n8534 = n8167 & ~n8422;
  assign n8535 = n8534 ^ n8169;
  assign n8536 = n8535 ^ n8532;
  assign n8537 = n8533 & ~n8536;
  assign n8538 = n8537 ^ n5625;
  assign n8539 = n8538 ^ n8439;
  assign n8540 = ~n8440 & n8539;
  assign n8541 = n8540 ^ n5363;
  assign n8542 = n8541 ^ n8436;
  assign n8543 = n8437 & ~n8542;
  assign n8544 = n8543 ^ n5108;
  assign n8545 = n8544 ^ n4851;
  assign n8546 = n8185 & ~n8422;
  assign n8547 = n8546 ^ n8187;
  assign n8548 = n8547 ^ n8544;
  assign n8549 = n8545 & n8548;
  assign n8550 = n8549 ^ n4851;
  assign n8551 = n8550 ^ n4606;
  assign n8552 = n8191 & ~n8422;
  assign n8553 = n8552 ^ n8193;
  assign n8554 = n8553 ^ n8550;
  assign n8555 = n8551 & ~n8554;
  assign n8556 = n8555 ^ n4606;
  assign n8557 = n8556 ^ n4362;
  assign n8558 = n8197 & ~n8422;
  assign n8559 = n8558 ^ n8199;
  assign n8560 = n8559 ^ n8556;
  assign n8561 = n8557 & n8560;
  assign n8562 = n8561 ^ n4362;
  assign n8563 = n8562 ^ n4133;
  assign n8564 = n8202 ^ n4362;
  assign n8565 = ~n8422 & n8564;
  assign n8566 = n8565 ^ n8085;
  assign n8567 = n8566 ^ n8562;
  assign n8568 = n8563 & ~n8567;
  assign n8569 = n8568 ^ n4133;
  assign n8570 = n8569 ^ n3882;
  assign n8571 = n8202 ^ n8085;
  assign n8572 = n8564 & ~n8571;
  assign n8573 = n8572 ^ n4362;
  assign n8574 = n8573 ^ n4133;
  assign n8575 = ~n8422 & n8574;
  assign n8576 = n8575 ^ n8088;
  assign n8577 = n8576 ^ n8569;
  assign n8578 = n8570 & n8577;
  assign n8579 = n8578 ^ n3882;
  assign n8580 = n8579 ^ n3634;
  assign n8581 = ~n8210 & ~n8422;
  assign n8582 = n8581 ^ n8212;
  assign n8583 = n8582 ^ n8579;
  assign n8584 = ~n8580 & ~n8583;
  assign n8585 = n8584 ^ n3634;
  assign n8586 = n8585 ^ n3397;
  assign n8587 = ~n8216 & ~n8422;
  assign n8588 = n8587 ^ n8219;
  assign n8589 = n8588 ^ n8585;
  assign n8590 = ~n8586 & ~n8589;
  assign n8591 = n8590 ^ n3397;
  assign n8592 = n8591 ^ n3177;
  assign n8593 = ~n8223 & ~n8422;
  assign n8594 = n8593 ^ n8226;
  assign n8595 = n8594 ^ n8591;
  assign n8596 = n8592 & ~n8595;
  assign n8597 = n8596 ^ n3177;
  assign n8598 = n8597 ^ n8433;
  assign n8599 = ~n8434 & n8598;
  assign n8600 = n8599 ^ n2980;
  assign n8601 = n8600 ^ n8430;
  assign n8602 = n8431 & ~n8601;
  assign n8603 = n8602 ^ n2782;
  assign n8604 = n8603 ^ n2583;
  assign n8605 = n8242 & ~n8422;
  assign n8606 = n8605 ^ n8244;
  assign n8607 = n8606 ^ n8603;
  assign n8608 = n8604 & n8607;
  assign n8609 = n8608 ^ n2583;
  assign n8610 = n8609 ^ n8427;
  assign n8611 = n8428 & ~n8610;
  assign n8612 = n8611 ^ n2374;
  assign n8613 = n8612 ^ n8424;
  assign n8614 = n8425 & n8613;
  assign n8615 = n8614 ^ n2194;
  assign n8616 = n8615 ^ n2011;
  assign n8617 = ~n8290 & ~n8422;
  assign n8618 = n8617 ^ n8292;
  assign n8619 = n8618 ^ n8615;
  assign n8620 = ~n8616 & n8619;
  assign n8621 = n8620 ^ n2011;
  assign n8622 = n8621 ^ n1804;
  assign n8623 = ~n8296 & ~n8422;
  assign n8624 = n8623 ^ n8298;
  assign n8625 = n8624 ^ n8621;
  assign n8626 = n8622 & n8625;
  assign n8627 = n8626 ^ n1804;
  assign n8628 = n8627 ^ n1621;
  assign n8629 = n8302 & ~n8422;
  assign n8630 = n8629 ^ n8304;
  assign n8631 = n8630 ^ n8627;
  assign n8632 = n8628 & ~n8631;
  assign n8633 = n8632 ^ n1621;
  assign n8634 = n8633 ^ n1458;
  assign n8635 = n8308 & ~n8422;
  assign n8636 = n8635 ^ n8310;
  assign n8637 = n8636 ^ n8633;
  assign n8638 = n8634 & n8637;
  assign n8639 = n8638 ^ n1458;
  assign n8640 = n8639 ^ n1299;
  assign n8641 = n8314 & ~n8422;
  assign n8642 = n8641 ^ n8316;
  assign n8643 = n8642 ^ n8639;
  assign n8644 = n8640 & ~n8643;
  assign n8645 = n8644 ^ n1299;
  assign n8646 = n8645 ^ n1158;
  assign n8647 = n8320 & ~n8422;
  assign n8648 = n8647 ^ n8322;
  assign n8649 = n8648 ^ n8645;
  assign n8650 = n8646 & n8649;
  assign n8651 = n8650 ^ n1158;
  assign n8652 = n8651 ^ n1027;
  assign n8653 = n8326 & ~n8422;
  assign n8654 = n8653 ^ n8328;
  assign n8655 = n8654 ^ n8651;
  assign n8656 = n8652 & ~n8655;
  assign n8657 = n8656 ^ n1027;
  assign n8658 = n8657 ^ n905;
  assign n8659 = n8332 & ~n8422;
  assign n8660 = n8659 ^ n8334;
  assign n8661 = n8660 ^ n8657;
  assign n8662 = n8658 & n8661;
  assign n8663 = n8662 ^ n905;
  assign n8664 = n8663 ^ n803;
  assign n8665 = n8338 & ~n8422;
  assign n8666 = n8665 ^ n8340;
  assign n8667 = n8666 ^ n8663;
  assign n8668 = n8664 & ~n8667;
  assign n8669 = n8668 ^ n803;
  assign n8670 = n8669 ^ n707;
  assign n8671 = ~n8379 & ~n8422;
  assign n8672 = n8671 ^ n8381;
  assign n8673 = ~n132 & n8672;
  assign n8674 = n8351 & ~n8422;
  assign n8675 = n8674 ^ n8353;
  assign n8676 = n8675 ^ n436;
  assign n8677 = n8275 ^ n803;
  assign n8678 = n8343 ^ n8275;
  assign n8679 = n8677 & ~n8678;
  assign n8680 = n8679 ^ n803;
  assign n8681 = n8680 ^ n8272;
  assign n8682 = ~n8273 & ~n8681;
  assign n8683 = n8682 ^ n707;
  assign n8684 = n8683 ^ n608;
  assign n8685 = ~n8422 & ~n8684;
  assign n8686 = n8685 ^ n8269;
  assign n8687 = n8686 ^ n514;
  assign n8688 = n8343 ^ n803;
  assign n8689 = ~n8422 & n8688;
  assign n8690 = n8689 ^ n8275;
  assign n8691 = n8690 ^ n8669;
  assign n8692 = ~n8670 & ~n8691;
  assign n8693 = n8692 ^ n707;
  assign n8694 = n8693 ^ n608;
  assign n8695 = n8680 ^ n707;
  assign n8696 = ~n8422 & ~n8695;
  assign n8697 = n8696 ^ n8272;
  assign n8698 = n8697 ^ n8693;
  assign n8699 = ~n8694 & n8698;
  assign n8700 = n8699 ^ n608;
  assign n8701 = n8700 ^ n8686;
  assign n8702 = ~n8687 & n8701;
  assign n8703 = n8702 ^ n514;
  assign n8704 = n8703 ^ n8675;
  assign n8705 = n8676 & ~n8704;
  assign n8706 = n8705 ^ n436;
  assign n8707 = n8706 ^ n363;
  assign n8708 = n8357 & ~n8422;
  assign n8709 = n8708 ^ n8360;
  assign n8710 = n8709 ^ n8706;
  assign n8711 = n8707 & n8710;
  assign n8712 = n8711 ^ n363;
  assign n8713 = n8712 ^ n300;
  assign n8714 = n8363 ^ n363;
  assign n8715 = ~n8422 & n8714;
  assign n8716 = n8715 ^ n8266;
  assign n8717 = n8716 ^ n8712;
  assign n8718 = n8713 & ~n8717;
  assign n8719 = n8718 ^ n300;
  assign n8720 = n8719 ^ n243;
  assign n8721 = n8366 ^ n300;
  assign n8722 = ~n8422 & n8721;
  assign n8723 = n8722 ^ n8262;
  assign n8724 = n8723 ^ n8719;
  assign n8725 = n8720 & ~n8724;
  assign n8726 = n8725 ^ n243;
  assign n8727 = n8726 ^ n210;
  assign n8728 = n8369 ^ n243;
  assign n8729 = ~n8422 & n8728;
  assign n8730 = n8729 ^ n8259;
  assign n8731 = n8730 ^ n8726;
  assign n8732 = n8727 & ~n8731;
  assign n8733 = n8732 ^ n210;
  assign n8734 = n8733 ^ n147;
  assign n8735 = n8373 & ~n8422;
  assign n8736 = n8735 ^ n8375;
  assign n8737 = n8736 ^ n8733;
  assign n8738 = ~n8734 & n8737;
  assign n8739 = n8738 ^ n147;
  assign n8740 = ~n8673 & n8739;
  assign n8741 = n8385 & ~n8422;
  assign n8742 = n8741 ^ n8387;
  assign n8743 = ~n133 & n8742;
  assign n8744 = n132 & ~n8672;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8740 & n8745;
  assign n8747 = n8387 & ~n8421;
  assign n8748 = ~n8256 & ~n8747;
  assign n8749 = n8393 ^ n7863;
  assign n8750 = ~n8053 & ~n8749;
  assign n8751 = n8750 ^ n7863;
  assign n8752 = n8751 ^ n133;
  assign n8753 = n8752 ^ n8751;
  assign n8754 = ~n8384 & ~n8387;
  assign n8755 = ~n132 & n8754;
  assign n8756 = n8755 ^ n8751;
  assign n8757 = n8753 & n8756;
  assign n8758 = n8757 ^ n8751;
  assign n8759 = ~n8390 & ~n8758;
  assign n8760 = n8759 ^ n133;
  assign n8761 = n8748 & n8760;
  assign n8762 = ~n133 & ~n8390;
  assign n8763 = n8384 & n8387;
  assign n8764 = n1292 & n8421;
  assign n8765 = n8763 & n8764;
  assign n8766 = n8256 & ~n8765;
  assign n8767 = ~n8762 & n8766;
  assign n8768 = ~n8761 & ~n8767;
  assign n8769 = ~n8746 & n8768;
  assign n8770 = ~n8670 & ~n8769;
  assign n8771 = n8770 ^ n8690;
  assign n8772 = n8771 ^ n608;
  assign n8773 = n8664 & ~n8769;
  assign n8774 = n8773 ^ n8666;
  assign n8775 = n8774 ^ n707;
  assign n8776 = n8612 ^ n2194;
  assign n8777 = ~n8769 & ~n8776;
  assign n8778 = n8777 ^ n8424;
  assign n8779 = n8778 ^ n2011;
  assign n8780 = n8609 ^ n2374;
  assign n8781 = ~n8769 & n8780;
  assign n8782 = n8781 ^ n8427;
  assign n8783 = n8782 ^ n2194;
  assign n8784 = n8597 ^ n2980;
  assign n8785 = ~n8769 & n8784;
  assign n8786 = n8785 ^ n8433;
  assign n8787 = n8786 ^ n2782;
  assign n8788 = n8592 & ~n8769;
  assign n8789 = n8788 ^ n8594;
  assign n8790 = n8789 ^ n2980;
  assign n8791 = n8533 & ~n8769;
  assign n8792 = n8791 ^ n8535;
  assign n8793 = n8792 ^ n5363;
  assign n8794 = n8527 & ~n8769;
  assign n8795 = n8794 ^ n8529;
  assign n8796 = n8795 ^ n5625;
  assign n8797 = n8463 & ~n8769;
  assign n8798 = ~x38 & ~n8797;
  assign n8799 = ~x34 & ~x35;
  assign n8800 = n8463 & n8799;
  assign n8801 = n8422 & n8800;
  assign n8802 = n8801 ^ x37;
  assign n8803 = n8802 ^ n8801;
  assign n8804 = ~x36 & n8799;
  assign n8805 = n8422 & ~n8804;
  assign n8806 = n8805 ^ n8801;
  assign n8807 = n8806 ^ n8801;
  assign n8808 = n8803 & n8807;
  assign n8809 = n8808 ^ n8801;
  assign n8810 = ~n8769 & ~n8809;
  assign n8811 = n8810 ^ n8801;
  assign n8812 = n8798 & n8811;
  assign n8813 = ~n8769 & ~n8800;
  assign n8814 = x37 & ~n8804;
  assign n8815 = n8461 & ~n8814;
  assign n8816 = ~n8813 & n8815;
  assign n8817 = ~n8812 & ~n8816;
  assign n8818 = ~n8422 & n8769;
  assign n8819 = x37 & n8818;
  assign n8820 = n8798 & ~n8819;
  assign n8821 = n8804 ^ x38;
  assign n8822 = x37 & n8821;
  assign n8823 = n8822 ^ x38;
  assign n8824 = ~n8769 & n8823;
  assign n8825 = n8422 ^ x38;
  assign n8826 = n8804 ^ n8422;
  assign n8827 = n8826 ^ n8804;
  assign n8828 = n8804 ^ n8800;
  assign n8829 = n8827 & ~n8828;
  assign n8830 = n8829 ^ n8804;
  assign n8831 = ~n8825 & n8830;
  assign n8832 = n8831 ^ x38;
  assign n8833 = ~n8824 & ~n8832;
  assign n8834 = ~n8820 & n8833;
  assign n8835 = ~n8083 & ~n8834;
  assign n8836 = n8817 & ~n8835;
  assign n8837 = n8836 ^ n7777;
  assign n8839 = n8422 ^ n8083;
  assign n8840 = n8839 ^ n8422;
  assign n8841 = n8840 ^ n8839;
  assign n8842 = n8839 ^ n8463;
  assign n8843 = n8841 & n8842;
  assign n8844 = n8843 ^ n8839;
  assign n8845 = ~x38 & n8844;
  assign n8846 = n8845 ^ n8839;
  assign n8838 = ~x38 & ~n8422;
  assign n8847 = n8846 ^ n8838;
  assign n8848 = n8463 ^ n8083;
  assign n8849 = n8848 ^ n8846;
  assign n8850 = n8846 ^ n8769;
  assign n8851 = ~n8846 & n8850;
  assign n8852 = n8851 ^ n8846;
  assign n8853 = ~n8849 & ~n8852;
  assign n8854 = n8853 ^ n8851;
  assign n8855 = n8854 ^ n8846;
  assign n8856 = n8855 ^ n8769;
  assign n8857 = n8847 & n8856;
  assign n8858 = n8857 ^ n8838;
  assign n8859 = n8858 ^ x39;
  assign n8860 = n8859 ^ n8836;
  assign n8861 = n8837 & ~n8860;
  assign n8862 = n8861 ^ n7777;
  assign n8863 = n8862 ^ n7463;
  assign n8864 = n8471 & ~n8769;
  assign n8865 = n8864 ^ n8475;
  assign n8866 = n8865 ^ n8862;
  assign n8867 = n8863 & n8866;
  assign n8868 = n8867 ^ n7463;
  assign n8869 = n8868 ^ n7135;
  assign n8870 = n8479 & ~n8769;
  assign n8871 = n8870 ^ n8497;
  assign n8872 = n8871 ^ n8868;
  assign n8873 = n8869 & ~n8872;
  assign n8874 = n8873 ^ n7135;
  assign n8875 = n8874 ^ n6802;
  assign n8876 = n8500 ^ n7135;
  assign n8877 = ~n8769 & n8876;
  assign n8878 = n8877 ^ n8459;
  assign n8879 = n8878 ^ n8874;
  assign n8880 = n8875 & ~n8879;
  assign n8881 = n8880 ^ n6802;
  assign n8882 = n8881 ^ n6479;
  assign n8883 = n8513 ^ n6802;
  assign n8884 = ~n8769 & n8883;
  assign n8885 = n8884 ^ n8507;
  assign n8886 = n8885 ^ n8881;
  assign n8887 = n8882 & ~n8886;
  assign n8888 = n8887 ^ n6479;
  assign n8889 = n8888 ^ n6181;
  assign n8890 = n8513 ^ n8507;
  assign n8891 = n8883 & ~n8890;
  assign n8892 = n8891 ^ n6802;
  assign n8893 = n8892 ^ n6479;
  assign n8894 = ~n8769 & n8893;
  assign n8895 = n8894 ^ n8443;
  assign n8896 = n8895 ^ n8888;
  assign n8897 = n8889 & n8896;
  assign n8898 = n8897 ^ n6181;
  assign n8899 = n8898 ^ n5905;
  assign n8900 = n8521 & ~n8769;
  assign n8901 = n8900 ^ n8523;
  assign n8902 = n8901 ^ n8898;
  assign n8903 = n8899 & ~n8902;
  assign n8904 = n8903 ^ n5905;
  assign n8905 = n8904 ^ n8795;
  assign n8906 = ~n8796 & n8905;
  assign n8907 = n8906 ^ n5625;
  assign n8908 = n8907 ^ n8792;
  assign n8909 = n8793 & ~n8908;
  assign n8910 = n8909 ^ n5363;
  assign n8911 = n8910 ^ n5108;
  assign n8912 = n8538 ^ n5363;
  assign n8913 = ~n8769 & n8912;
  assign n8914 = n8913 ^ n8439;
  assign n8915 = n8914 ^ n8910;
  assign n8916 = n8911 & n8915;
  assign n8917 = n8916 ^ n5108;
  assign n8918 = n8917 ^ n4851;
  assign n8919 = n8541 ^ n5108;
  assign n8920 = ~n8769 & n8919;
  assign n8921 = n8920 ^ n8436;
  assign n8922 = n8921 ^ n8917;
  assign n8923 = n8918 & ~n8922;
  assign n8924 = n8923 ^ n4851;
  assign n8925 = n8924 ^ n4606;
  assign n8926 = n8545 & ~n8769;
  assign n8927 = n8926 ^ n8547;
  assign n8928 = n8927 ^ n8924;
  assign n8929 = n8925 & n8928;
  assign n8930 = n8929 ^ n4606;
  assign n8931 = n8930 ^ n4362;
  assign n8932 = n8551 & ~n8769;
  assign n8933 = n8932 ^ n8553;
  assign n8934 = n8933 ^ n8930;
  assign n8935 = n8931 & ~n8934;
  assign n8936 = n8935 ^ n4362;
  assign n8937 = n8936 ^ n4133;
  assign n8938 = n8557 & ~n8769;
  assign n8939 = n8938 ^ n8559;
  assign n8940 = n8939 ^ n8936;
  assign n8941 = n8937 & n8940;
  assign n8942 = n8941 ^ n4133;
  assign n8943 = n8942 ^ n3882;
  assign n8944 = n8563 & ~n8769;
  assign n8945 = n8944 ^ n8566;
  assign n8946 = n8945 ^ n8942;
  assign n8947 = n8943 & ~n8946;
  assign n8948 = n8947 ^ n3882;
  assign n8949 = n8948 ^ n3634;
  assign n8950 = n8570 & ~n8769;
  assign n8951 = n8950 ^ n8576;
  assign n8952 = n8951 ^ n8948;
  assign n8953 = ~n8949 & n8952;
  assign n8954 = n8953 ^ n3634;
  assign n8955 = n8954 ^ n3397;
  assign n8956 = ~n8580 & ~n8769;
  assign n8957 = n8956 ^ n8582;
  assign n8958 = n8957 ^ n8954;
  assign n8959 = ~n8955 & n8958;
  assign n8960 = n8959 ^ n3397;
  assign n8961 = n8960 ^ n3177;
  assign n8962 = ~n8586 & ~n8769;
  assign n8963 = n8962 ^ n8588;
  assign n8964 = n8963 ^ n8960;
  assign n8965 = n8961 & n8964;
  assign n8966 = n8965 ^ n3177;
  assign n8967 = n8966 ^ n8789;
  assign n8968 = n8790 & ~n8967;
  assign n8969 = n8968 ^ n2980;
  assign n8970 = n8969 ^ n8786;
  assign n8971 = ~n8787 & n8970;
  assign n8972 = n8971 ^ n2782;
  assign n8973 = n8972 ^ n2583;
  assign n8974 = n8600 ^ n2782;
  assign n8975 = ~n8769 & n8974;
  assign n8976 = n8975 ^ n8430;
  assign n8977 = n8976 ^ n8972;
  assign n8978 = n8973 & ~n8977;
  assign n8979 = n8978 ^ n2583;
  assign n8980 = n8979 ^ n2374;
  assign n8981 = n8604 & ~n8769;
  assign n8982 = n8981 ^ n8606;
  assign n8983 = n8982 ^ n8979;
  assign n8984 = n8980 & n8983;
  assign n8985 = n8984 ^ n2374;
  assign n8986 = n8985 ^ n8782;
  assign n8987 = ~n8783 & ~n8986;
  assign n8988 = n8987 ^ n2194;
  assign n8989 = n8988 ^ n8778;
  assign n8990 = ~n8779 & ~n8989;
  assign n8991 = n8990 ^ n2011;
  assign n8992 = n8991 ^ n1804;
  assign n8993 = ~n8616 & ~n8769;
  assign n8994 = n8993 ^ n8618;
  assign n8995 = n8994 ^ n8991;
  assign n8996 = n8992 & ~n8995;
  assign n8997 = n8996 ^ n1804;
  assign n8998 = n8997 ^ n1621;
  assign n8999 = n8622 & ~n8769;
  assign n9000 = n8999 ^ n8624;
  assign n9001 = n9000 ^ n8997;
  assign n9002 = n8998 & n9001;
  assign n9003 = n9002 ^ n1621;
  assign n9004 = n9003 ^ n1458;
  assign n9005 = n8628 & ~n8769;
  assign n9006 = n9005 ^ n8630;
  assign n9007 = n9006 ^ n9003;
  assign n9008 = n9004 & ~n9007;
  assign n9009 = n9008 ^ n1458;
  assign n9010 = n9009 ^ n1299;
  assign n9011 = n8634 & ~n8769;
  assign n9012 = n9011 ^ n8636;
  assign n9013 = n9012 ^ n9009;
  assign n9014 = n9010 & n9013;
  assign n9015 = n9014 ^ n1299;
  assign n9016 = n9015 ^ n1158;
  assign n9017 = n8640 & ~n8769;
  assign n9018 = n9017 ^ n8642;
  assign n9019 = n9018 ^ n9015;
  assign n9020 = n9016 & ~n9019;
  assign n9021 = n9020 ^ n1158;
  assign n9022 = n9021 ^ n1027;
  assign n9023 = n8646 & ~n8769;
  assign n9024 = n9023 ^ n8648;
  assign n9025 = n9024 ^ n9021;
  assign n9026 = n9022 & n9025;
  assign n9027 = n9026 ^ n1027;
  assign n9028 = n9027 ^ n905;
  assign n9029 = n8652 & ~n8769;
  assign n9030 = n9029 ^ n8654;
  assign n9031 = n9030 ^ n9027;
  assign n9032 = n9028 & ~n9031;
  assign n9033 = n9032 ^ n905;
  assign n9034 = n9033 ^ n803;
  assign n9035 = n8658 & ~n8769;
  assign n9036 = n9035 ^ n8660;
  assign n9037 = n9036 ^ n9033;
  assign n9038 = n9034 & n9037;
  assign n9039 = n9038 ^ n803;
  assign n9040 = n9039 ^ n8774;
  assign n9041 = ~n8775 & ~n9040;
  assign n9042 = n9041 ^ n707;
  assign n9043 = n9042 ^ n8771;
  assign n9044 = n8772 & n9043;
  assign n9045 = n9044 ^ n608;
  assign n9046 = n9045 ^ n514;
  assign n9047 = ~n8694 & ~n8769;
  assign n9048 = n9047 ^ n8697;
  assign n9049 = n9048 ^ n9045;
  assign n9050 = n9046 & ~n9049;
  assign n9051 = n9050 ^ n514;
  assign n9052 = n9051 ^ n436;
  assign n9053 = n8700 ^ n514;
  assign n9054 = ~n8769 & n9053;
  assign n9055 = n9054 ^ n8686;
  assign n9056 = n9055 ^ n9051;
  assign n9057 = n9052 & n9056;
  assign n9058 = n9057 ^ n436;
  assign n9059 = n9058 ^ n363;
  assign n9060 = n8703 ^ n436;
  assign n9061 = ~n8769 & n9060;
  assign n9062 = n9061 ^ n8675;
  assign n9063 = n9062 ^ n9058;
  assign n9064 = n9059 & ~n9063;
  assign n9065 = n9064 ^ n363;
  assign n9066 = n9065 ^ n300;
  assign n9067 = n8707 & ~n8769;
  assign n9068 = n9067 ^ n8709;
  assign n9069 = n9068 ^ n9065;
  assign n9070 = n9066 & n9069;
  assign n9071 = n9070 ^ n300;
  assign n9072 = n9071 ^ n243;
  assign n9073 = n8713 & ~n8769;
  assign n9074 = n9073 ^ n8716;
  assign n9075 = n9074 ^ n9071;
  assign n9076 = n9072 & ~n9075;
  assign n9077 = n9076 ^ n243;
  assign n9078 = n9077 ^ n210;
  assign n9079 = n8720 & ~n8769;
  assign n9080 = n9079 ^ n8723;
  assign n9081 = n9080 ^ n9077;
  assign n9082 = n9078 & ~n9081;
  assign n9083 = n9082 ^ n210;
  assign n9084 = n9083 ^ n147;
  assign n9085 = n8727 & ~n8769;
  assign n9086 = n9085 ^ n8730;
  assign n9087 = n9086 ^ n9083;
  assign n9088 = ~n9084 & ~n9087;
  assign n9089 = n9088 ^ n147;
  assign n9090 = n132 & n9089;
  assign n9091 = ~n8734 & ~n8769;
  assign n9092 = n9091 ^ n8736;
  assign n9093 = ~n9090 & ~n9092;
  assign n9094 = ~n132 & ~n9089;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = n8739 ^ n132;
  assign n9097 = ~n8769 & n9096;
  assign n9098 = n9097 ^ n8672;
  assign n9099 = ~n133 & ~n9098;
  assign n9100 = ~n9095 & ~n9099;
  assign n9101 = n8739 & ~n8742;
  assign n9102 = ~n8768 & ~n9101;
  assign n9103 = n133 & ~n8672;
  assign n9104 = ~n9102 & n9103;
  assign n9105 = n8672 & ~n8739;
  assign n9106 = n132 & ~n8743;
  assign n9107 = ~n9105 & n9106;
  assign n9108 = ~n9104 & n9107;
  assign n9109 = n8743 & ~n8768;
  assign n9110 = ~n8744 & n9109;
  assign n9111 = ~n8740 & n9110;
  assign n9112 = n8742 ^ n133;
  assign n9113 = n9112 ^ n8742;
  assign n9114 = n129 & ~n8768;
  assign n9115 = n9114 ^ n8742;
  assign n9116 = n9113 & ~n9115;
  assign n9117 = n9116 ^ n8742;
  assign n9118 = ~n8672 & ~n9117;
  assign n9119 = n8739 & n9118;
  assign n9120 = ~n9111 & ~n9119;
  assign n9121 = n8742 ^ n8672;
  assign n9122 = ~n132 & ~n8739;
  assign n9123 = n9122 ^ n8672;
  assign n9124 = ~n9121 & n9123;
  assign n9125 = n9124 ^ n8672;
  assign n9126 = n133 & n9125;
  assign n9127 = n9120 & ~n9126;
  assign n9128 = ~n9108 & n9127;
  assign n9129 = ~n9100 & n9128;
  assign n9130 = n8969 ^ n2782;
  assign n9131 = ~n9129 & n9130;
  assign n9132 = n9131 ^ n8786;
  assign n9133 = ~n2583 & n9132;
  assign n9134 = n8973 & ~n9129;
  assign n9135 = n9134 ^ n8976;
  assign n9136 = ~n2374 & ~n9135;
  assign n9137 = ~n9133 & ~n9136;
  assign n9138 = n8937 & ~n9129;
  assign n9139 = n9138 ^ n8939;
  assign n9140 = ~n3882 & n9139;
  assign n9141 = n8943 & ~n9129;
  assign n9142 = n9141 ^ n8945;
  assign n9143 = n3634 & ~n9142;
  assign n9144 = ~n9140 & ~n9143;
  assign n9145 = n8931 & ~n9129;
  assign n9146 = n9145 ^ n8933;
  assign n9147 = n9146 ^ n4133;
  assign n9148 = n8925 & ~n9129;
  assign n9149 = n9148 ^ n8927;
  assign n9150 = n9149 ^ n4362;
  assign n9151 = n8907 ^ n5363;
  assign n9152 = ~n9129 & n9151;
  assign n9153 = n9152 ^ n8792;
  assign n9154 = n9153 ^ n5108;
  assign n9155 = n8904 ^ n5625;
  assign n9156 = ~n9129 & n9155;
  assign n9157 = n9156 ^ n8795;
  assign n9158 = n9157 ^ n5363;
  assign n9159 = ~x32 & ~x33;
  assign n9160 = ~n8769 & n9159;
  assign n9161 = ~x34 & n9160;
  assign n9162 = n9129 ^ x35;
  assign n9163 = x34 & n8769;
  assign n9164 = n8769 & ~n9159;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = n9165 ^ x34;
  assign n9167 = n9166 ^ n9165;
  assign n9168 = n9165 ^ n9129;
  assign n9169 = n9168 ^ n9165;
  assign n9170 = n9167 & ~n9169;
  assign n9171 = n9170 ^ n9165;
  assign n9172 = ~n9162 & n9171;
  assign n9173 = n9172 ^ n9165;
  assign n9174 = ~n9161 & ~n9173;
  assign n9175 = n9174 ^ n8422;
  assign n9176 = n8799 ^ n8769;
  assign n9177 = ~n9129 & ~n9176;
  assign n9178 = n9177 ^ n8769;
  assign n9179 = n9178 ^ x36;
  assign n9180 = n9179 ^ n9174;
  assign n9181 = n9175 & n9180;
  assign n9182 = n9181 ^ n8422;
  assign n9183 = n9182 ^ n8083;
  assign n9185 = x36 & n8422;
  assign n9186 = n9185 ^ n8826;
  assign n9187 = ~n8769 & ~n9186;
  assign n9188 = n9187 ^ n8826;
  assign n9184 = ~x36 & ~n8769;
  assign n9189 = n9188 ^ n9184;
  assign n9190 = n8799 ^ n8422;
  assign n9191 = n9190 ^ n9188;
  assign n9192 = n9188 ^ n9129;
  assign n9193 = n9188 & ~n9192;
  assign n9194 = n9193 ^ n9188;
  assign n9195 = n9191 & n9194;
  assign n9196 = n9195 ^ n9193;
  assign n9197 = n9196 ^ n9188;
  assign n9198 = n9197 ^ n9129;
  assign n9199 = ~n9189 & ~n9198;
  assign n9200 = n9199 ^ n9184;
  assign n9201 = n9200 ^ x37;
  assign n9202 = n9201 ^ n9182;
  assign n9203 = n9183 & ~n9202;
  assign n9204 = n9203 ^ n8083;
  assign n9205 = n9204 ^ n7777;
  assign n9215 = ~n8797 & ~n8818;
  assign n9216 = n9215 ^ x38;
  assign n9206 = x36 & ~x37;
  assign n9207 = ~n8769 & n9206;
  assign n9208 = n8769 ^ x37;
  assign n9209 = n9208 ^ n8804;
  assign n9210 = ~n8826 & n9209;
  assign n9211 = n9210 ^ n8804;
  assign n9212 = ~n9207 & ~n9211;
  assign n9213 = n9212 ^ n8083;
  assign n9214 = ~n9129 & n9213;
  assign n9217 = n9216 ^ n9214;
  assign n9218 = n9217 ^ n9204;
  assign n9219 = n9205 & n9218;
  assign n9220 = n9219 ^ n7777;
  assign n9221 = n9220 ^ n7463;
  assign n9222 = n8859 ^ n7777;
  assign n9223 = n9222 ^ n8817;
  assign n9224 = n9223 ^ n8834;
  assign n9225 = n9224 ^ n9222;
  assign n9226 = n8834 ^ n8083;
  assign n9227 = n9226 ^ n8083;
  assign n9228 = n9222 ^ n8083;
  assign n9229 = n9227 & ~n9228;
  assign n9230 = n9229 ^ n8083;
  assign n9231 = n9225 & ~n9230;
  assign n9232 = n9231 ^ n9223;
  assign n9233 = n9232 ^ n8859;
  assign n9234 = ~n9129 & n9233;
  assign n9235 = n9234 ^ n8859;
  assign n9236 = n9235 ^ n9220;
  assign n9237 = n9221 & ~n9236;
  assign n9238 = n9237 ^ n7463;
  assign n9239 = n9238 ^ n7135;
  assign n9240 = n8863 & ~n9129;
  assign n9241 = n9240 ^ n8865;
  assign n9242 = n9241 ^ n9238;
  assign n9243 = n9239 & n9242;
  assign n9244 = n9243 ^ n7135;
  assign n9245 = n9244 ^ n6802;
  assign n9246 = n8869 & ~n9129;
  assign n9247 = n9246 ^ n8871;
  assign n9248 = n9247 ^ n9244;
  assign n9249 = n9245 & ~n9248;
  assign n9250 = n9249 ^ n6802;
  assign n9251 = n9250 ^ n6479;
  assign n9252 = n8875 & ~n9129;
  assign n9253 = n9252 ^ n8878;
  assign n9254 = n9253 ^ n9250;
  assign n9255 = n9251 & ~n9254;
  assign n9256 = n9255 ^ n6479;
  assign n9257 = n9256 ^ n6181;
  assign n9258 = n8882 & ~n9129;
  assign n9259 = n9258 ^ n8885;
  assign n9260 = n9259 ^ n9256;
  assign n9261 = n9257 & ~n9260;
  assign n9262 = n9261 ^ n6181;
  assign n9263 = n9262 ^ n5905;
  assign n9264 = n8889 & ~n9129;
  assign n9265 = n9264 ^ n8895;
  assign n9266 = n9265 ^ n9262;
  assign n9267 = n9263 & n9266;
  assign n9268 = n9267 ^ n5905;
  assign n9269 = n9268 ^ n5625;
  assign n9270 = n8899 & ~n9129;
  assign n9271 = n9270 ^ n8901;
  assign n9272 = n9271 ^ n9268;
  assign n9273 = n9269 & ~n9272;
  assign n9274 = n9273 ^ n5625;
  assign n9275 = n9274 ^ n9157;
  assign n9276 = ~n9158 & n9275;
  assign n9277 = n9276 ^ n5363;
  assign n9278 = n9277 ^ n9153;
  assign n9279 = n9154 & ~n9278;
  assign n9280 = n9279 ^ n5108;
  assign n9281 = n9280 ^ n4851;
  assign n9282 = n8911 & ~n9129;
  assign n9283 = n9282 ^ n8914;
  assign n9284 = n9283 ^ n9280;
  assign n9285 = n9281 & n9284;
  assign n9286 = n9285 ^ n4851;
  assign n9287 = n9286 ^ n4606;
  assign n9288 = n8918 & ~n9129;
  assign n9289 = n9288 ^ n8921;
  assign n9290 = n9289 ^ n9286;
  assign n9291 = n9287 & ~n9290;
  assign n9292 = n9291 ^ n4606;
  assign n9293 = n9292 ^ n9149;
  assign n9294 = ~n9150 & n9293;
  assign n9295 = n9294 ^ n4362;
  assign n9296 = n9295 ^ n9146;
  assign n9297 = n9147 & ~n9296;
  assign n9298 = n9297 ^ n4133;
  assign n9299 = n9144 & n9298;
  assign n9300 = ~n8949 & ~n9129;
  assign n9301 = n9300 ^ n8951;
  assign n9302 = n3397 & ~n9301;
  assign n9303 = ~n8955 & ~n9129;
  assign n9304 = n9303 ^ n8957;
  assign n9305 = n3177 & n9304;
  assign n9306 = ~n9302 & ~n9305;
  assign n9307 = n9142 ^ n3634;
  assign n9308 = n3882 & ~n9139;
  assign n9309 = n9308 ^ n9142;
  assign n9310 = ~n9307 & ~n9309;
  assign n9311 = n9310 ^ n3634;
  assign n9312 = n9306 & n9311;
  assign n9313 = ~n9299 & n9312;
  assign n9314 = n9304 ^ n3177;
  assign n9315 = ~n3397 & n9301;
  assign n9316 = n9315 ^ n9304;
  assign n9317 = n9314 & n9316;
  assign n9318 = n9317 ^ n3177;
  assign n9319 = ~n9313 & n9318;
  assign n9320 = n9319 ^ n2980;
  assign n9321 = n8961 & ~n9129;
  assign n9322 = n9321 ^ n8963;
  assign n9323 = n9322 ^ n9319;
  assign n9324 = n9320 & n9323;
  assign n9325 = n9324 ^ n2980;
  assign n9326 = n9325 ^ n2782;
  assign n9327 = n8966 ^ n2980;
  assign n9328 = ~n9129 & n9327;
  assign n9329 = n9328 ^ n8789;
  assign n9330 = n9329 ^ n9325;
  assign n9331 = n9326 & ~n9330;
  assign n9332 = n9331 ^ n2782;
  assign n9333 = n9137 & n9332;
  assign n9334 = n9135 ^ n2374;
  assign n9335 = n2583 & ~n9132;
  assign n9336 = n9335 ^ n9135;
  assign n9337 = n9334 & ~n9336;
  assign n9338 = n9337 ^ n2374;
  assign n9339 = ~n9333 & ~n9338;
  assign n9340 = n9339 ^ n2194;
  assign n9341 = n8980 & ~n9129;
  assign n9342 = n9341 ^ n8982;
  assign n9343 = n9342 ^ n9339;
  assign n9344 = n9340 & ~n9343;
  assign n9345 = n9344 ^ n2194;
  assign n9346 = n9345 ^ n2011;
  assign n9347 = n8985 ^ n2194;
  assign n9348 = ~n9129 & ~n9347;
  assign n9349 = n9348 ^ n8782;
  assign n9350 = n9349 ^ n9345;
  assign n9351 = ~n9346 & n9350;
  assign n9352 = n9351 ^ n2011;
  assign n9353 = n9352 ^ n1804;
  assign n9354 = n8988 ^ n2011;
  assign n9355 = ~n9129 & ~n9354;
  assign n9356 = n9355 ^ n8778;
  assign n9357 = n9356 ^ n9352;
  assign n9358 = n9353 & n9357;
  assign n9359 = n9358 ^ n1804;
  assign n9360 = n9359 ^ n1621;
  assign n9361 = n8992 & ~n9129;
  assign n9362 = n9361 ^ n8994;
  assign n9363 = n9362 ^ n9359;
  assign n9364 = n9360 & ~n9363;
  assign n9365 = n9364 ^ n1621;
  assign n9366 = n9365 ^ n1458;
  assign n9367 = n8998 & ~n9129;
  assign n9368 = n9367 ^ n9000;
  assign n9369 = n9368 ^ n9365;
  assign n9370 = n9366 & n9369;
  assign n9371 = n9370 ^ n1458;
  assign n9372 = n9371 ^ n1299;
  assign n9373 = n9004 & ~n9129;
  assign n9374 = n9373 ^ n9006;
  assign n9375 = n9374 ^ n9371;
  assign n9376 = n9372 & ~n9375;
  assign n9377 = n9376 ^ n1299;
  assign n9378 = n9377 ^ n1158;
  assign n9379 = n9010 & ~n9129;
  assign n9380 = n9379 ^ n9012;
  assign n9381 = n9380 ^ n9377;
  assign n9382 = n9378 & n9381;
  assign n9383 = n9382 ^ n1158;
  assign n9384 = n9383 ^ n1027;
  assign n9385 = n9016 & ~n9129;
  assign n9386 = n9385 ^ n9018;
  assign n9387 = n9386 ^ n9383;
  assign n9388 = n9384 & ~n9387;
  assign n9389 = n9388 ^ n1027;
  assign n9390 = n9389 ^ n905;
  assign n9391 = n9022 & ~n9129;
  assign n9392 = n9391 ^ n9024;
  assign n9393 = n9392 ^ n9389;
  assign n9394 = n9390 & n9393;
  assign n9395 = n9394 ^ n905;
  assign n9396 = n9395 ^ n803;
  assign n9397 = n9028 & ~n9129;
  assign n9398 = n9397 ^ n9030;
  assign n9399 = n9398 ^ n9395;
  assign n9400 = n9396 & ~n9399;
  assign n9401 = n9400 ^ n803;
  assign n9402 = n9401 ^ n707;
  assign n9403 = n9034 & ~n9129;
  assign n9404 = n9403 ^ n9036;
  assign n9405 = n9404 ^ n9401;
  assign n9406 = ~n9402 & n9405;
  assign n9407 = n9406 ^ n707;
  assign n9408 = n9407 ^ n608;
  assign n9409 = n9039 ^ n707;
  assign n9410 = ~n9129 & ~n9409;
  assign n9411 = n9410 ^ n8774;
  assign n9412 = n9411 ^ n9407;
  assign n9413 = ~n9408 & n9412;
  assign n9414 = n9413 ^ n608;
  assign n9415 = n9414 ^ n514;
  assign n9416 = n9042 ^ n608;
  assign n9417 = ~n9129 & ~n9416;
  assign n9418 = n9417 ^ n8771;
  assign n9419 = n9418 ^ n9414;
  assign n9420 = n9415 & ~n9419;
  assign n9421 = n9420 ^ n514;
  assign n9422 = n9421 ^ n436;
  assign n9423 = n9046 & ~n9129;
  assign n9424 = n9423 ^ n9048;
  assign n9425 = n9424 ^ n9421;
  assign n9426 = n9422 & ~n9425;
  assign n9427 = n9426 ^ n436;
  assign n9428 = n9427 ^ n363;
  assign n9429 = n9052 & ~n9129;
  assign n9430 = n9429 ^ n9055;
  assign n9431 = n9430 ^ n9427;
  assign n9432 = n9428 & n9431;
  assign n9433 = n9432 ^ n363;
  assign n9434 = n9433 ^ n300;
  assign n9435 = n9078 & ~n9129;
  assign n9436 = n9435 ^ n9080;
  assign n9437 = n9066 & ~n9129;
  assign n9438 = n9437 ^ n9068;
  assign n9439 = n9438 ^ n243;
  assign n9440 = n9059 & ~n9129;
  assign n9441 = n9440 ^ n9062;
  assign n9442 = n9441 ^ n9433;
  assign n9443 = n9434 & ~n9442;
  assign n9444 = n9443 ^ n300;
  assign n9445 = n9444 ^ n9438;
  assign n9446 = ~n9439 & n9445;
  assign n9447 = n9446 ^ n243;
  assign n9448 = n9447 ^ n210;
  assign n9449 = n9072 & ~n9129;
  assign n9450 = n9449 ^ n9074;
  assign n9451 = n9450 ^ n9447;
  assign n9452 = n9448 & ~n9451;
  assign n9453 = n9452 ^ n210;
  assign n9454 = ~n9436 & ~n9453;
  assign n9455 = n1973 & ~n9454;
  assign n9456 = ~n9084 & ~n9129;
  assign n9457 = n9456 ^ n9086;
  assign n9458 = n9457 ^ n9436;
  assign n9459 = n9457 ^ n132;
  assign n9460 = n9459 ^ n132;
  assign n9461 = ~n182 & n9460;
  assign n9462 = n9461 ^ n132;
  assign n9463 = n9458 & n9462;
  assign n9464 = n9463 ^ n9436;
  assign n9465 = n9453 & n9464;
  assign n9466 = n9436 ^ n147;
  assign n9467 = ~n147 & ~n182;
  assign n9468 = n9467 ^ n147;
  assign n9469 = ~n9466 & ~n9468;
  assign n9470 = n9469 ^ n9467;
  assign n9471 = n9470 ^ n147;
  assign n9472 = n9471 ^ n132;
  assign n9473 = n9457 & ~n9472;
  assign n9474 = n9473 ^ n9457;
  assign n9475 = ~n9465 & ~n9474;
  assign n9476 = ~n9455 & n9475;
  assign n9477 = n9089 ^ n132;
  assign n9478 = ~n9129 & n9477;
  assign n9479 = n9478 ^ n9092;
  assign n9480 = ~n133 & n9479;
  assign n9481 = ~n9476 & ~n9480;
  assign n9483 = ~n9098 & n9128;
  assign n9484 = n9483 ^ n9094;
  assign n9485 = n9093 & ~n9484;
  assign n9482 = n9098 ^ n9094;
  assign n9486 = n9485 ^ n9482;
  assign n9487 = ~n133 & ~n9486;
  assign n9488 = n9092 & n9483;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = n9092 ^ n9089;
  assign n9491 = ~n132 & ~n9490;
  assign n9492 = n133 & ~n9491;
  assign n9493 = n9089 & n9092;
  assign n9494 = ~n9128 & n9493;
  assign n9495 = n9494 ^ n9098;
  assign n9496 = n9495 ^ n9494;
  assign n9497 = n9494 ^ n9095;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = n9498 ^ n9494;
  assign n9500 = n9492 & n9499;
  assign n9501 = n9489 & ~n9500;
  assign n9502 = ~n9481 & ~n9501;
  assign n9503 = n9434 & ~n9502;
  assign n9504 = n9503 ^ n9441;
  assign n9505 = n9504 ^ n243;
  assign n9506 = n9428 & ~n9502;
  assign n9507 = n9506 ^ n9430;
  assign n9508 = n9507 ^ n300;
  assign n9509 = n9422 & ~n9502;
  assign n9510 = n9509 ^ n9424;
  assign n9511 = n9510 ^ n363;
  assign n9512 = ~n9408 & ~n9502;
  assign n9513 = n9512 ^ n9411;
  assign n9514 = n9513 ^ n514;
  assign n9515 = ~n9402 & ~n9502;
  assign n9516 = n9515 ^ n9404;
  assign n9517 = n9516 ^ n608;
  assign n9518 = ~n9299 & n9311;
  assign n9519 = n9518 ^ n3397;
  assign n9520 = ~n9502 & ~n9519;
  assign n9521 = n9520 ^ n9301;
  assign n9522 = n9521 ^ n3177;
  assign n9523 = n9298 ^ n3882;
  assign n9524 = n9298 ^ n9139;
  assign n9525 = n9523 & n9524;
  assign n9526 = n9525 ^ n3882;
  assign n9527 = n9526 ^ n3634;
  assign n9528 = ~n9502 & ~n9527;
  assign n9529 = n9528 ^ n9142;
  assign n9530 = n9529 ^ n3397;
  assign n9531 = n9281 & ~n9502;
  assign n9532 = n9531 ^ n9283;
  assign n9533 = n9532 ^ n4606;
  assign n9534 = n9277 ^ n5108;
  assign n9535 = ~n9502 & n9534;
  assign n9536 = n9535 ^ n9153;
  assign n9537 = n9536 ^ n4851;
  assign n9538 = n9221 & ~n9502;
  assign n9539 = n9538 ^ n9235;
  assign n9540 = n9539 ^ n7135;
  assign n9541 = n9205 & ~n9502;
  assign n9542 = n9541 ^ n9217;
  assign n9543 = n9542 ^ n7463;
  assign n9544 = ~x30 & ~x31;
  assign n9545 = ~x32 & n9544;
  assign n9546 = n9129 & ~n9545;
  assign n9547 = n9502 ^ x33;
  assign n9548 = ~n9546 & n9547;
  assign n9550 = ~n9129 & n9544;
  assign n9549 = ~x33 & ~n9502;
  assign n9551 = n9550 ^ n9549;
  assign n9552 = ~x32 & n9551;
  assign n9553 = n9552 ^ n9549;
  assign n9554 = ~n9548 & ~n9553;
  assign n9555 = n9554 ^ n8769;
  assign n9556 = n9159 ^ n9129;
  assign n9557 = ~n9502 & ~n9556;
  assign n9558 = n9557 ^ n9129;
  assign n9559 = n9558 ^ x34;
  assign n9560 = n9559 ^ n9554;
  assign n9561 = n9555 & n9560;
  assign n9562 = n9561 ^ n8769;
  assign n9563 = n9562 ^ n8422;
  assign n9565 = n9163 ^ n9161;
  assign n9566 = n9565 ^ n9163;
  assign n9567 = n9165 ^ n9163;
  assign n9568 = n9567 ^ n9163;
  assign n9569 = ~n9566 & n9568;
  assign n9570 = n9569 ^ n9163;
  assign n9571 = n9129 & n9570;
  assign n9572 = n9571 ^ n9163;
  assign n9564 = ~x34 & ~n9129;
  assign n9573 = n9572 ^ n9564;
  assign n9574 = n9159 ^ n8769;
  assign n9575 = n9574 ^ n9572;
  assign n9576 = n9572 ^ n9502;
  assign n9577 = ~n9572 & n9576;
  assign n9578 = n9577 ^ n9572;
  assign n9579 = ~n9575 & ~n9578;
  assign n9580 = n9579 ^ n9577;
  assign n9581 = n9580 ^ n9572;
  assign n9582 = n9581 ^ n9502;
  assign n9583 = n9573 & n9582;
  assign n9584 = n9583 ^ n9564;
  assign n9585 = n9584 ^ x35;
  assign n9586 = n9585 ^ n9562;
  assign n9587 = n9563 & ~n9586;
  assign n9588 = n9587 ^ n8422;
  assign n9589 = n9588 ^ n8083;
  assign n9590 = n9175 & ~n9502;
  assign n9591 = n9590 ^ n9179;
  assign n9592 = n9591 ^ n9588;
  assign n9593 = n9589 & n9592;
  assign n9594 = n9593 ^ n8083;
  assign n9595 = n9594 ^ n7777;
  assign n9596 = n9183 & ~n9502;
  assign n9597 = n9596 ^ n9201;
  assign n9598 = n9597 ^ n9594;
  assign n9599 = n9595 & ~n9598;
  assign n9600 = n9599 ^ n7777;
  assign n9601 = n9600 ^ n9542;
  assign n9602 = ~n9543 & n9601;
  assign n9603 = n9602 ^ n7463;
  assign n9604 = n9603 ^ n9539;
  assign n9605 = n9540 & ~n9604;
  assign n9606 = n9605 ^ n7135;
  assign n9607 = n9606 ^ n6802;
  assign n9608 = n9239 & ~n9502;
  assign n9609 = n9608 ^ n9241;
  assign n9610 = n9609 ^ n9606;
  assign n9611 = n9607 & n9610;
  assign n9612 = n9611 ^ n6802;
  assign n9613 = n9612 ^ n6479;
  assign n9614 = n9245 & ~n9502;
  assign n9615 = n9614 ^ n9247;
  assign n9616 = n9615 ^ n9612;
  assign n9617 = n9613 & ~n9616;
  assign n9618 = n9617 ^ n6479;
  assign n9619 = n9618 ^ n6181;
  assign n9620 = n9251 & ~n9502;
  assign n9621 = n9620 ^ n9253;
  assign n9622 = n9621 ^ n9618;
  assign n9623 = n9619 & ~n9622;
  assign n9624 = n9623 ^ n6181;
  assign n9625 = n9624 ^ n5905;
  assign n9626 = n9257 & ~n9502;
  assign n9627 = n9626 ^ n9259;
  assign n9628 = n9627 ^ n9624;
  assign n9629 = n9625 & ~n9628;
  assign n9630 = n9629 ^ n5905;
  assign n9631 = n9630 ^ n5625;
  assign n9632 = n9263 & ~n9502;
  assign n9633 = n9632 ^ n9265;
  assign n9634 = n9633 ^ n9630;
  assign n9635 = n9631 & n9634;
  assign n9636 = n9635 ^ n5625;
  assign n9637 = n9636 ^ n5363;
  assign n9638 = n9269 & ~n9502;
  assign n9639 = n9638 ^ n9271;
  assign n9640 = n9639 ^ n9636;
  assign n9641 = n9637 & ~n9640;
  assign n9642 = n9641 ^ n5363;
  assign n9643 = n9642 ^ n5108;
  assign n9644 = n9274 ^ n5363;
  assign n9645 = ~n9502 & n9644;
  assign n9646 = n9645 ^ n9157;
  assign n9647 = n9646 ^ n9642;
  assign n9648 = n9643 & n9647;
  assign n9649 = n9648 ^ n5108;
  assign n9650 = n9649 ^ n9536;
  assign n9651 = n9537 & ~n9650;
  assign n9652 = n9651 ^ n4851;
  assign n9653 = n9652 ^ n9532;
  assign n9654 = ~n9533 & n9653;
  assign n9655 = n9654 ^ n4606;
  assign n9656 = n9655 ^ n4362;
  assign n9657 = n9287 & ~n9502;
  assign n9658 = n9657 ^ n9289;
  assign n9659 = n9658 ^ n9655;
  assign n9660 = n9656 & ~n9659;
  assign n9661 = n9660 ^ n4362;
  assign n9662 = n9661 ^ n4133;
  assign n9663 = n9292 ^ n4362;
  assign n9664 = ~n9502 & n9663;
  assign n9665 = n9664 ^ n9149;
  assign n9666 = n9665 ^ n9661;
  assign n9667 = n9662 & n9666;
  assign n9668 = n9667 ^ n4133;
  assign n9669 = n9668 ^ n3882;
  assign n9670 = n9295 ^ n4133;
  assign n9671 = ~n9502 & n9670;
  assign n9672 = n9671 ^ n9146;
  assign n9673 = n9672 ^ n9668;
  assign n9674 = n9669 & ~n9673;
  assign n9675 = n9674 ^ n3882;
  assign n9676 = n9675 ^ n3634;
  assign n9677 = ~n9502 & n9523;
  assign n9678 = n9677 ^ n9139;
  assign n9679 = n9678 ^ n9675;
  assign n9680 = ~n9676 & n9679;
  assign n9681 = n9680 ^ n3634;
  assign n9682 = n9681 ^ n9529;
  assign n9683 = n9530 & n9682;
  assign n9684 = n9683 ^ n3397;
  assign n9685 = n9684 ^ n9521;
  assign n9686 = ~n9522 & n9685;
  assign n9687 = n9686 ^ n3177;
  assign n9688 = n9687 ^ n2980;
  assign n9689 = n9301 ^ n3397;
  assign n9690 = n9518 ^ n9301;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n9691 ^ n3397;
  assign n9693 = n9692 ^ n3177;
  assign n9694 = ~n9502 & n9693;
  assign n9695 = n9694 ^ n9304;
  assign n9696 = n9695 ^ n9687;
  assign n9697 = n9688 & ~n9696;
  assign n9698 = n9697 ^ n2980;
  assign n9699 = n9698 ^ n2782;
  assign n9700 = n9320 & ~n9502;
  assign n9701 = n9700 ^ n9322;
  assign n9702 = n9701 ^ n9698;
  assign n9703 = n9699 & n9702;
  assign n9704 = n9703 ^ n2782;
  assign n9705 = n9704 ^ n2583;
  assign n9706 = n9326 & ~n9502;
  assign n9707 = n9706 ^ n9329;
  assign n9708 = n9707 ^ n9704;
  assign n9709 = n9705 & ~n9708;
  assign n9710 = n9709 ^ n2583;
  assign n9711 = n9710 ^ n2374;
  assign n9712 = n9332 ^ n2583;
  assign n9713 = ~n9502 & n9712;
  assign n9714 = n9713 ^ n9132;
  assign n9715 = n9714 ^ n9710;
  assign n9716 = n9711 & n9715;
  assign n9717 = n9716 ^ n2374;
  assign n9718 = n9717 ^ n2194;
  assign n9719 = n9332 ^ n9132;
  assign n9720 = n9712 & n9719;
  assign n9721 = n9720 ^ n2583;
  assign n9722 = n9721 ^ n2374;
  assign n9723 = ~n9502 & n9722;
  assign n9724 = n9723 ^ n9135;
  assign n9725 = n9724 ^ n9717;
  assign n9726 = ~n9718 & ~n9725;
  assign n9727 = n9726 ^ n2194;
  assign n9728 = n9727 ^ n2011;
  assign n9729 = n9340 & ~n9502;
  assign n9730 = n9729 ^ n9342;
  assign n9731 = n9730 ^ n9727;
  assign n9732 = ~n9728 & ~n9731;
  assign n9733 = n9732 ^ n2011;
  assign n9734 = n9733 ^ n1804;
  assign n9735 = ~n9346 & ~n9502;
  assign n9736 = n9735 ^ n9349;
  assign n9737 = n9736 ^ n9733;
  assign n9738 = n9734 & ~n9737;
  assign n9739 = n9738 ^ n1804;
  assign n9740 = n9739 ^ n1621;
  assign n9741 = n9353 & ~n9502;
  assign n9742 = n9741 ^ n9356;
  assign n9743 = n9742 ^ n9739;
  assign n9744 = n9740 & n9743;
  assign n9745 = n9744 ^ n1621;
  assign n9746 = n9745 ^ n1458;
  assign n9747 = n9360 & ~n9502;
  assign n9748 = n9747 ^ n9362;
  assign n9749 = n9748 ^ n9745;
  assign n9750 = n9746 & ~n9749;
  assign n9751 = n9750 ^ n1458;
  assign n9752 = n9751 ^ n1299;
  assign n9753 = n9366 & ~n9502;
  assign n9754 = n9753 ^ n9368;
  assign n9755 = n9754 ^ n9751;
  assign n9756 = n9752 & n9755;
  assign n9757 = n9756 ^ n1299;
  assign n9758 = n9757 ^ n1158;
  assign n9759 = n9372 & ~n9502;
  assign n9760 = n9759 ^ n9374;
  assign n9761 = n9760 ^ n9757;
  assign n9762 = n9758 & ~n9761;
  assign n9763 = n9762 ^ n1158;
  assign n9764 = n9763 ^ n1027;
  assign n9765 = n9378 & ~n9502;
  assign n9766 = n9765 ^ n9380;
  assign n9767 = n9766 ^ n9763;
  assign n9768 = n9764 & n9767;
  assign n9769 = n9768 ^ n1027;
  assign n9770 = n9769 ^ n905;
  assign n9771 = n9384 & ~n9502;
  assign n9772 = n9771 ^ n9386;
  assign n9773 = n9772 ^ n9769;
  assign n9774 = n9770 & ~n9773;
  assign n9775 = n9774 ^ n905;
  assign n9776 = n9775 ^ n803;
  assign n9777 = n9390 & ~n9502;
  assign n9778 = n9777 ^ n9392;
  assign n9779 = n9778 ^ n9775;
  assign n9780 = n9776 & n9779;
  assign n9781 = n9780 ^ n803;
  assign n9782 = n9781 ^ n707;
  assign n9783 = n9396 & ~n9502;
  assign n9784 = n9783 ^ n9398;
  assign n9785 = n9784 ^ n9781;
  assign n9786 = ~n9782 & ~n9785;
  assign n9787 = n9786 ^ n707;
  assign n9788 = n9787 ^ n9516;
  assign n9789 = ~n9517 & ~n9788;
  assign n9790 = n9789 ^ n608;
  assign n9791 = n9790 ^ n9513;
  assign n9792 = n9514 & ~n9791;
  assign n9793 = n9792 ^ n514;
  assign n9794 = n9793 ^ n436;
  assign n9795 = n9415 & ~n9502;
  assign n9796 = n9795 ^ n9418;
  assign n9797 = n9796 ^ n9793;
  assign n9798 = n9794 & ~n9797;
  assign n9799 = n9798 ^ n436;
  assign n9800 = n9799 ^ n9510;
  assign n9801 = n9511 & ~n9800;
  assign n9802 = n9801 ^ n363;
  assign n9803 = n9802 ^ n9507;
  assign n9804 = ~n9508 & n9803;
  assign n9805 = n9804 ^ n300;
  assign n9806 = n9805 ^ n9504;
  assign n9807 = n9505 & ~n9806;
  assign n9808 = n9807 ^ n243;
  assign n9809 = n9808 ^ n210;
  assign n9810 = n9444 ^ n243;
  assign n9811 = ~n9502 & n9810;
  assign n9812 = n9811 ^ n9438;
  assign n9813 = n9812 ^ n9808;
  assign n9814 = n9809 & n9813;
  assign n9815 = n9814 ^ n210;
  assign n9816 = n9815 ^ n147;
  assign n9817 = n9448 & ~n9502;
  assign n9818 = n9817 ^ n9450;
  assign n9819 = n9818 ^ n9815;
  assign n9820 = ~n9816 & ~n9819;
  assign n9821 = n9820 ^ n147;
  assign n9822 = n132 & n9821;
  assign n9823 = n9453 ^ n147;
  assign n9824 = ~n9502 & ~n9823;
  assign n9825 = n9824 ^ n9436;
  assign n9826 = ~n9822 & n9825;
  assign n9827 = ~n132 & ~n9821;
  assign n9828 = ~n9826 & ~n9827;
  assign n9829 = n9453 ^ n9436;
  assign n9830 = ~n9823 & ~n9829;
  assign n9831 = n9830 ^ n147;
  assign n9832 = n9831 ^ n132;
  assign n9833 = ~n9502 & n9832;
  assign n9834 = n9833 ^ n9457;
  assign n9835 = ~n133 & ~n9834;
  assign n9836 = ~n9828 & ~n9835;
  assign n9837 = ~n132 & ~n9831;
  assign n9838 = n9501 ^ n9479;
  assign n9839 = n133 & ~n9838;
  assign n9840 = n9839 ^ n9479;
  assign n9841 = ~n9837 & n9840;
  assign n9842 = n9479 ^ n132;
  assign n9843 = n9831 ^ n9479;
  assign n9844 = n9842 & n9843;
  assign n9845 = n133 & n9844;
  assign n9846 = ~n9841 & ~n9845;
  assign n9847 = ~n9457 & ~n9846;
  assign n9848 = n1287 & n9457;
  assign n9849 = n9831 & n9848;
  assign n9850 = ~n133 & ~n9489;
  assign n9851 = n9479 & ~n9850;
  assign n9852 = ~n9849 & n9851;
  assign n9853 = n9831 ^ n133;
  assign n9854 = n9831 ^ n9457;
  assign n9855 = ~n9831 & ~n9832;
  assign n9856 = n9855 ^ n9831;
  assign n9857 = n9854 & ~n9856;
  assign n9858 = n9857 ^ n9855;
  assign n9859 = n9858 ^ n9831;
  assign n9860 = n9859 ^ n132;
  assign n9861 = n9853 & ~n9860;
  assign n9862 = n9852 & ~n9861;
  assign n9863 = ~n133 & ~n9476;
  assign n9864 = ~n9479 & ~n9863;
  assign n9865 = ~n9862 & ~n9864;
  assign n9866 = ~n9847 & ~n9865;
  assign n9867 = ~n9836 & ~n9866;
  assign n9868 = ~n9816 & ~n9867;
  assign n9869 = n9868 ^ n9818;
  assign n9870 = n132 & ~n9869;
  assign n9871 = n9752 & ~n9867;
  assign n9872 = n9871 ^ n9754;
  assign n9873 = n9872 ^ n1158;
  assign n9874 = n9746 & ~n9867;
  assign n9875 = n9874 ^ n9748;
  assign n9876 = n9875 ^ n1299;
  assign n9877 = n9669 & ~n9867;
  assign n9878 = n9877 ^ n9672;
  assign n9879 = n9878 ^ n3634;
  assign n9880 = n9662 & ~n9867;
  assign n9881 = n9880 ^ n9665;
  assign n9882 = n9881 ^ n3882;
  assign n9883 = ~x28 & ~x29;
  assign n9884 = ~n9502 & n9883;
  assign n9885 = ~x30 & n9884;
  assign n9892 = n9867 ^ n9544;
  assign n9893 = n9892 ^ x31;
  assign n9886 = n9502 & n9883;
  assign n9887 = ~x30 & n9886;
  assign n9888 = n9887 ^ n9502;
  assign n9894 = n9888 ^ x31;
  assign n9895 = n9894 ^ n9544;
  assign n9896 = ~n9893 & n9895;
  assign n9898 = n9896 ^ n9885;
  assign n9889 = n9888 ^ n9544;
  assign n9890 = n9889 ^ n9544;
  assign n9891 = ~n9889 & ~n9890;
  assign n9899 = n9891 ^ n9889;
  assign n9900 = n9898 & ~n9899;
  assign n9897 = n9896 ^ n9891;
  assign n9901 = n9900 ^ n9897;
  assign n9902 = n9885 & n9901;
  assign n9903 = n9902 ^ n9896;
  assign n9904 = n9903 ^ n9891;
  assign n9905 = n9904 ^ n9900;
  assign n9906 = n9905 ^ n9885;
  assign n9907 = n9906 ^ n9129;
  assign n9908 = n9544 ^ n9502;
  assign n9909 = ~n9867 & ~n9908;
  assign n9910 = n9909 ^ n9502;
  assign n9911 = n9910 ^ x32;
  assign n9912 = n9911 ^ n9906;
  assign n9913 = ~n9907 & ~n9912;
  assign n9914 = n9913 ^ n9129;
  assign n9915 = n9914 ^ n8769;
  assign n9917 = n9545 ^ n9129;
  assign n9918 = n9917 ^ x32;
  assign n9919 = n9918 ^ n9917;
  assign n9920 = n9917 ^ n9545;
  assign n9921 = n9919 & n9920;
  assign n9922 = n9921 ^ n9917;
  assign n9923 = ~n9502 & ~n9922;
  assign n9924 = n9923 ^ n9917;
  assign n9916 = ~x32 & ~n9502;
  assign n9925 = n9924 ^ n9916;
  assign n9926 = n9544 ^ n9129;
  assign n9927 = n9926 ^ n9924;
  assign n9928 = n9924 ^ n9867;
  assign n9929 = n9924 & ~n9928;
  assign n9930 = n9929 ^ n9924;
  assign n9931 = n9927 & n9930;
  assign n9932 = n9931 ^ n9929;
  assign n9933 = n9932 ^ n9924;
  assign n9934 = n9933 ^ n9867;
  assign n9935 = ~n9925 & ~n9934;
  assign n9936 = n9935 ^ n9916;
  assign n9937 = n9936 ^ x33;
  assign n9938 = n9937 ^ n9914;
  assign n9939 = n9915 & ~n9938;
  assign n9940 = n9939 ^ n8769;
  assign n9941 = n9940 ^ n8422;
  assign n9942 = n9555 & ~n9867;
  assign n9943 = n9942 ^ n9559;
  assign n9944 = n9943 ^ n9940;
  assign n9945 = n9941 & n9944;
  assign n9946 = n9945 ^ n8422;
  assign n9947 = n9946 ^ n8083;
  assign n9948 = n9563 & ~n9867;
  assign n9949 = n9948 ^ n9585;
  assign n9950 = n9949 ^ n9946;
  assign n9951 = n9947 & ~n9950;
  assign n9952 = n9951 ^ n8083;
  assign n9953 = n9952 ^ n7777;
  assign n9954 = n9589 & ~n9867;
  assign n9955 = n9954 ^ n9591;
  assign n9956 = n9955 ^ n9952;
  assign n9957 = n9953 & n9956;
  assign n9958 = n9957 ^ n7777;
  assign n9959 = n9958 ^ n7463;
  assign n9960 = n9595 & ~n9867;
  assign n9961 = n9960 ^ n9597;
  assign n9962 = n9961 ^ n9958;
  assign n9963 = n9959 & ~n9962;
  assign n9964 = n9963 ^ n7463;
  assign n9965 = n9964 ^ n7135;
  assign n9966 = n9600 ^ n7463;
  assign n9967 = ~n9867 & n9966;
  assign n9968 = n9967 ^ n9542;
  assign n9969 = n9968 ^ n9964;
  assign n9970 = n9965 & n9969;
  assign n9971 = n9970 ^ n7135;
  assign n9972 = n9971 ^ n6802;
  assign n9973 = n9603 ^ n7135;
  assign n9974 = ~n9867 & n9973;
  assign n9975 = n9974 ^ n9539;
  assign n9976 = n9975 ^ n9971;
  assign n9977 = n9972 & ~n9976;
  assign n9978 = n9977 ^ n6802;
  assign n9979 = n9978 ^ n6479;
  assign n9980 = n9607 & ~n9867;
  assign n9981 = n9980 ^ n9609;
  assign n9982 = n9981 ^ n9978;
  assign n9983 = n9979 & n9982;
  assign n9984 = n9983 ^ n6479;
  assign n9985 = n9984 ^ n6181;
  assign n9986 = n9613 & ~n9867;
  assign n9987 = n9986 ^ n9615;
  assign n9988 = n9987 ^ n9984;
  assign n9989 = n9985 & ~n9988;
  assign n9990 = n9989 ^ n6181;
  assign n9991 = n9990 ^ n5905;
  assign n9992 = n9619 & ~n9867;
  assign n9993 = n9992 ^ n9621;
  assign n9994 = n9993 ^ n9990;
  assign n9995 = n9991 & ~n9994;
  assign n9996 = n9995 ^ n5905;
  assign n9997 = n9996 ^ n5625;
  assign n9998 = n9625 & ~n9867;
  assign n9999 = n9998 ^ n9627;
  assign n10000 = n9999 ^ n9996;
  assign n10001 = n9997 & ~n10000;
  assign n10002 = n10001 ^ n5625;
  assign n10003 = n10002 ^ n5363;
  assign n10004 = n9631 & ~n9867;
  assign n10005 = n10004 ^ n9633;
  assign n10006 = n10005 ^ n10002;
  assign n10007 = n10003 & n10006;
  assign n10008 = n10007 ^ n5363;
  assign n10009 = n10008 ^ n5108;
  assign n10010 = n9637 & ~n9867;
  assign n10011 = n10010 ^ n9639;
  assign n10012 = n10011 ^ n10008;
  assign n10013 = n10009 & ~n10012;
  assign n10014 = n10013 ^ n5108;
  assign n10015 = n10014 ^ n4851;
  assign n10016 = n9643 & ~n9867;
  assign n10017 = n10016 ^ n9646;
  assign n10018 = n10017 ^ n10014;
  assign n10019 = n10015 & n10018;
  assign n10020 = n10019 ^ n4851;
  assign n10021 = n10020 ^ n4606;
  assign n10022 = n9649 ^ n4851;
  assign n10023 = ~n9867 & n10022;
  assign n10024 = n10023 ^ n9536;
  assign n10025 = n10024 ^ n10020;
  assign n10026 = n10021 & ~n10025;
  assign n10027 = n10026 ^ n4606;
  assign n10028 = n10027 ^ n4362;
  assign n10029 = n9652 ^ n4606;
  assign n10030 = ~n9867 & n10029;
  assign n10031 = n10030 ^ n9532;
  assign n10032 = n10031 ^ n10027;
  assign n10033 = n10028 & n10032;
  assign n10034 = n10033 ^ n4362;
  assign n10035 = n10034 ^ n4133;
  assign n10036 = n9656 & ~n9867;
  assign n10037 = n10036 ^ n9658;
  assign n10038 = n10037 ^ n10034;
  assign n10039 = n10035 & ~n10038;
  assign n10040 = n10039 ^ n4133;
  assign n10041 = n10040 ^ n9881;
  assign n10042 = ~n9882 & n10041;
  assign n10043 = n10042 ^ n3882;
  assign n10044 = n10043 ^ n9878;
  assign n10045 = ~n9879 & ~n10044;
  assign n10046 = n10045 ^ n3634;
  assign n10047 = n10046 ^ n3397;
  assign n10048 = ~n9676 & ~n9867;
  assign n10049 = n10048 ^ n9678;
  assign n10050 = n10049 ^ n10046;
  assign n10051 = ~n10047 & ~n10050;
  assign n10052 = n10051 ^ n3397;
  assign n10053 = n10052 ^ n3177;
  assign n10054 = n9681 ^ n3397;
  assign n10055 = ~n9867 & ~n10054;
  assign n10056 = n10055 ^ n9529;
  assign n10057 = n10056 ^ n10052;
  assign n10058 = n10053 & ~n10057;
  assign n10059 = n10058 ^ n3177;
  assign n10060 = n10059 ^ n2980;
  assign n10061 = n9684 ^ n3177;
  assign n10062 = ~n9867 & n10061;
  assign n10063 = n10062 ^ n9521;
  assign n10064 = n10063 ^ n10059;
  assign n10065 = n10060 & n10064;
  assign n10066 = n10065 ^ n2980;
  assign n10067 = n10066 ^ n2782;
  assign n10068 = n9688 & ~n9867;
  assign n10069 = n10068 ^ n9695;
  assign n10070 = n10069 ^ n10066;
  assign n10071 = n10067 & ~n10070;
  assign n10072 = n10071 ^ n2782;
  assign n10073 = n10072 ^ n2583;
  assign n10074 = n9699 & ~n9867;
  assign n10075 = n10074 ^ n9701;
  assign n10076 = n10075 ^ n10072;
  assign n10077 = n10073 & n10076;
  assign n10078 = n10077 ^ n2583;
  assign n10079 = n10078 ^ n2374;
  assign n10080 = n9705 & ~n9867;
  assign n10081 = n10080 ^ n9707;
  assign n10082 = n10081 ^ n10078;
  assign n10083 = n10079 & ~n10082;
  assign n10084 = n10083 ^ n2374;
  assign n10085 = n10084 ^ n2194;
  assign n10086 = n9711 & ~n9867;
  assign n10087 = n10086 ^ n9714;
  assign n10088 = n10087 ^ n10084;
  assign n10089 = ~n10085 & n10088;
  assign n10090 = n10089 ^ n2194;
  assign n10091 = n10090 ^ n2011;
  assign n10092 = ~n9718 & ~n9867;
  assign n10093 = n10092 ^ n9724;
  assign n10094 = n10093 ^ n10090;
  assign n10095 = ~n10091 & n10094;
  assign n10096 = n10095 ^ n2011;
  assign n10097 = n10096 ^ n1804;
  assign n10098 = ~n9728 & ~n9867;
  assign n10099 = n10098 ^ n9730;
  assign n10100 = n10099 ^ n10096;
  assign n10101 = n10097 & n10100;
  assign n10102 = n10101 ^ n1804;
  assign n10103 = n10102 ^ n1621;
  assign n10104 = n9734 & ~n9867;
  assign n10105 = n10104 ^ n9736;
  assign n10106 = n10105 ^ n10102;
  assign n10107 = n10103 & ~n10106;
  assign n10108 = n10107 ^ n1621;
  assign n10109 = n10108 ^ n1458;
  assign n10110 = n9740 & ~n9867;
  assign n10111 = n10110 ^ n9742;
  assign n10112 = n10111 ^ n10108;
  assign n10113 = n10109 & n10112;
  assign n10114 = n10113 ^ n1458;
  assign n10115 = n10114 ^ n9875;
  assign n10116 = n9876 & ~n10115;
  assign n10117 = n10116 ^ n1299;
  assign n10118 = n10117 ^ n9872;
  assign n10119 = ~n9873 & n10118;
  assign n10120 = n10119 ^ n1158;
  assign n10121 = n10120 ^ n1027;
  assign n10122 = n9758 & ~n9867;
  assign n10123 = n10122 ^ n9760;
  assign n10124 = n10123 ^ n10120;
  assign n10125 = n10121 & ~n10124;
  assign n10126 = n10125 ^ n1027;
  assign n10127 = n10126 ^ n905;
  assign n10128 = n9764 & ~n9867;
  assign n10129 = n10128 ^ n9766;
  assign n10130 = n10129 ^ n10126;
  assign n10131 = n10127 & n10130;
  assign n10132 = n10131 ^ n905;
  assign n10133 = n10132 ^ n803;
  assign n10134 = n9770 & ~n9867;
  assign n10135 = n10134 ^ n9772;
  assign n10136 = n10135 ^ n10132;
  assign n10137 = n10133 & ~n10136;
  assign n10138 = n10137 ^ n803;
  assign n10139 = n10138 ^ n707;
  assign n10140 = n9776 & ~n9867;
  assign n10141 = n10140 ^ n9778;
  assign n10142 = n10141 ^ n10138;
  assign n10143 = ~n10139 & n10142;
  assign n10144 = n10143 ^ n707;
  assign n10145 = n10144 ^ n608;
  assign n10146 = ~n9782 & ~n9867;
  assign n10147 = n10146 ^ n9784;
  assign n10148 = n10147 ^ n10144;
  assign n10149 = ~n10145 & n10148;
  assign n10150 = n10149 ^ n608;
  assign n10151 = n10150 ^ n514;
  assign n10152 = n9787 ^ n608;
  assign n10153 = ~n9867 & ~n10152;
  assign n10154 = n10153 ^ n9516;
  assign n10155 = n10154 ^ n10150;
  assign n10156 = n10151 & n10155;
  assign n10157 = n10156 ^ n514;
  assign n10158 = n10157 ^ n436;
  assign n10159 = n9790 ^ n514;
  assign n10160 = ~n9867 & n10159;
  assign n10161 = n10160 ^ n9513;
  assign n10162 = n10161 ^ n10157;
  assign n10163 = n10158 & ~n10162;
  assign n10164 = n10163 ^ n436;
  assign n10165 = n10164 ^ n363;
  assign n10166 = n9794 & ~n9867;
  assign n10167 = n10166 ^ n9796;
  assign n10168 = n10167 ^ n10164;
  assign n10169 = n10165 & ~n10168;
  assign n10170 = n10169 ^ n363;
  assign n10171 = n10170 ^ n300;
  assign n10172 = n9799 ^ n363;
  assign n10173 = ~n9867 & n10172;
  assign n10174 = n10173 ^ n9510;
  assign n10175 = n10174 ^ n10170;
  assign n10176 = n10171 & ~n10175;
  assign n10177 = n10176 ^ n300;
  assign n10178 = n10177 ^ n243;
  assign n10179 = n9802 ^ n300;
  assign n10180 = ~n9867 & n10179;
  assign n10181 = n10180 ^ n9507;
  assign n10182 = n10181 ^ n10177;
  assign n10183 = n10178 & n10182;
  assign n10184 = n10183 ^ n243;
  assign n10185 = n10184 ^ n210;
  assign n10186 = n9805 ^ n243;
  assign n10187 = ~n9867 & n10186;
  assign n10188 = n10187 ^ n9504;
  assign n10189 = n10188 ^ n10184;
  assign n10190 = n10185 & ~n10189;
  assign n10191 = n10190 ^ n210;
  assign n10192 = n10191 ^ n147;
  assign n10193 = n9809 & ~n9867;
  assign n10194 = n10193 ^ n9812;
  assign n10195 = n10194 ^ n10191;
  assign n10196 = ~n10192 & n10195;
  assign n10197 = n10196 ^ n147;
  assign n10198 = ~n9870 & ~n10197;
  assign n10199 = ~n132 & n9869;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = n9821 ^ n132;
  assign n10202 = ~n9867 & n10201;
  assign n10203 = n10202 ^ n9825;
  assign n10204 = ~n133 & ~n10203;
  assign n10205 = ~n10200 & ~n10204;
  assign n10206 = ~n9827 & n9866;
  assign n10207 = ~n9825 & ~n10206;
  assign n10208 = n133 & ~n9834;
  assign n10209 = ~n10207 & n10208;
  assign n10210 = n9826 & ~n9827;
  assign n10211 = n10209 & ~n10210;
  assign n10216 = n9835 & n9866;
  assign n10212 = n1292 & ~n9825;
  assign n10213 = n9866 & n10212;
  assign n10214 = n9821 & n10213;
  assign n10215 = n9834 & ~n10214;
  assign n10217 = n10216 ^ n10215;
  assign n10218 = n10216 ^ n133;
  assign n10219 = n10216 ^ n9828;
  assign n10220 = ~n10216 & n10219;
  assign n10221 = n10220 ^ n10216;
  assign n10222 = ~n10218 & ~n10221;
  assign n10223 = n10222 ^ n10220;
  assign n10224 = n10223 ^ n10216;
  assign n10225 = n10224 ^ n9828;
  assign n10226 = n10217 & n10225;
  assign n10227 = n10226 ^ n10215;
  assign n10228 = ~n10211 & ~n10227;
  assign n10229 = ~n10205 & n10228;
  assign n10230 = n10117 ^ n1158;
  assign n10231 = ~n10229 & n10230;
  assign n10232 = n10231 ^ n9872;
  assign n10233 = n10232 ^ n1027;
  assign n10234 = n10114 ^ n1299;
  assign n10235 = ~n10229 & n10234;
  assign n10236 = n10235 ^ n9875;
  assign n10237 = n10236 ^ n1158;
  assign n10238 = n10109 & ~n10229;
  assign n10239 = n10238 ^ n10111;
  assign n10240 = n10239 ^ n1299;
  assign n10241 = n10103 & ~n10229;
  assign n10242 = n10241 ^ n10105;
  assign n10243 = n10242 ^ n1458;
  assign n10244 = n10073 & ~n10229;
  assign n10245 = n10244 ^ n10075;
  assign n10246 = n10245 ^ n2374;
  assign n10247 = n10067 & ~n10229;
  assign n10248 = n10247 ^ n10069;
  assign n10249 = n10248 ^ n2583;
  assign n10250 = x28 & n9867;
  assign n10251 = ~x26 & ~x27;
  assign n10252 = n9867 & ~n10251;
  assign n10253 = ~n10250 & ~n10252;
  assign n10254 = n10229 ^ x29;
  assign n10255 = n10253 & n10254;
  assign n10257 = ~n9867 & n10251;
  assign n10256 = ~x29 & ~n10229;
  assign n10258 = n10257 ^ n10256;
  assign n10259 = ~x28 & n10258;
  assign n10260 = n10259 ^ n10256;
  assign n10261 = ~n10255 & ~n10260;
  assign n10262 = n10261 ^ n9502;
  assign n10263 = n9883 ^ n9867;
  assign n10264 = ~n10229 & ~n10263;
  assign n10265 = n10264 ^ n9867;
  assign n10266 = n10265 ^ x30;
  assign n10267 = n10266 ^ n10261;
  assign n10268 = n10262 & n10267;
  assign n10269 = n10268 ^ n9502;
  assign n10270 = n10269 ^ n9129;
  assign n10272 = n9867 ^ n9502;
  assign n10273 = n10272 ^ n9867;
  assign n10274 = n10273 ^ n10272;
  assign n10275 = n10272 ^ n9883;
  assign n10276 = n10274 & n10275;
  assign n10277 = n10276 ^ n10272;
  assign n10278 = ~x30 & n10277;
  assign n10279 = n10278 ^ n10272;
  assign n10271 = ~x30 & ~n9867;
  assign n10280 = n10279 ^ n10271;
  assign n10281 = n9883 ^ n9502;
  assign n10282 = n10281 ^ n10279;
  assign n10283 = n10279 ^ n10229;
  assign n10284 = ~n10279 & n10283;
  assign n10285 = n10284 ^ n10279;
  assign n10286 = ~n10282 & ~n10285;
  assign n10287 = n10286 ^ n10284;
  assign n10288 = n10287 ^ n10279;
  assign n10289 = n10288 ^ n10229;
  assign n10290 = n10280 & n10289;
  assign n10291 = n10290 ^ n10271;
  assign n10292 = n10291 ^ x31;
  assign n10293 = n10292 ^ n10269;
  assign n10294 = n10270 & ~n10293;
  assign n10295 = n10294 ^ n9129;
  assign n10296 = n10295 ^ n8769;
  assign n10297 = ~n9907 & ~n10229;
  assign n10298 = n10297 ^ n9911;
  assign n10299 = n10298 ^ n10295;
  assign n10300 = n10296 & n10299;
  assign n10301 = n10300 ^ n8769;
  assign n10302 = n10301 ^ n8422;
  assign n10303 = n9915 & ~n10229;
  assign n10304 = n10303 ^ n9937;
  assign n10305 = n10304 ^ n10301;
  assign n10306 = n10302 & ~n10305;
  assign n10307 = n10306 ^ n8422;
  assign n10308 = n10307 ^ n8083;
  assign n10309 = n9941 & ~n10229;
  assign n10310 = n10309 ^ n9943;
  assign n10311 = n10310 ^ n10307;
  assign n10312 = n10308 & n10311;
  assign n10313 = n10312 ^ n8083;
  assign n10314 = n10313 ^ n7777;
  assign n10315 = n9947 & ~n10229;
  assign n10316 = n10315 ^ n9949;
  assign n10317 = n10316 ^ n10313;
  assign n10318 = n10314 & ~n10317;
  assign n10319 = n10318 ^ n7777;
  assign n10320 = n10319 ^ n7463;
  assign n10321 = n9953 & ~n10229;
  assign n10322 = n10321 ^ n9955;
  assign n10323 = n10322 ^ n10319;
  assign n10324 = n10320 & n10323;
  assign n10325 = n10324 ^ n7463;
  assign n10326 = n10325 ^ n7135;
  assign n10327 = n9959 & ~n10229;
  assign n10328 = n10327 ^ n9961;
  assign n10329 = n10328 ^ n10325;
  assign n10330 = n10326 & ~n10329;
  assign n10331 = n10330 ^ n7135;
  assign n10332 = n10331 ^ n6802;
  assign n10333 = n9965 & ~n10229;
  assign n10334 = n10333 ^ n9968;
  assign n10335 = n10334 ^ n10331;
  assign n10336 = n10332 & n10335;
  assign n10337 = n10336 ^ n6802;
  assign n10338 = n10337 ^ n6479;
  assign n10339 = n9972 & ~n10229;
  assign n10340 = n10339 ^ n9975;
  assign n10341 = n10340 ^ n10337;
  assign n10342 = n10338 & ~n10341;
  assign n10343 = n10342 ^ n6479;
  assign n10344 = n10343 ^ n6181;
  assign n10345 = n9979 & ~n10229;
  assign n10346 = n10345 ^ n9981;
  assign n10347 = n10346 ^ n10343;
  assign n10348 = n10344 & n10347;
  assign n10349 = n10348 ^ n6181;
  assign n10350 = n10349 ^ n5905;
  assign n10351 = n9985 & ~n10229;
  assign n10352 = n10351 ^ n9987;
  assign n10353 = n10352 ^ n10349;
  assign n10354 = n10350 & ~n10353;
  assign n10355 = n10354 ^ n5905;
  assign n10356 = n10355 ^ n5625;
  assign n10357 = n9991 & ~n10229;
  assign n10358 = n10357 ^ n9993;
  assign n10359 = n10358 ^ n10355;
  assign n10360 = n10356 & ~n10359;
  assign n10361 = n10360 ^ n5625;
  assign n10362 = n10361 ^ n5363;
  assign n10363 = n9997 & ~n10229;
  assign n10364 = n10363 ^ n9999;
  assign n10365 = n10364 ^ n10361;
  assign n10366 = n10362 & ~n10365;
  assign n10367 = n10366 ^ n5363;
  assign n10368 = n10367 ^ n5108;
  assign n10369 = n10003 & ~n10229;
  assign n10370 = n10369 ^ n10005;
  assign n10371 = n10370 ^ n10367;
  assign n10372 = n10368 & n10371;
  assign n10373 = n10372 ^ n5108;
  assign n10374 = n10373 ^ n4851;
  assign n10375 = n10009 & ~n10229;
  assign n10376 = n10375 ^ n10011;
  assign n10377 = n10376 ^ n10373;
  assign n10378 = n10374 & ~n10377;
  assign n10379 = n10378 ^ n4851;
  assign n10380 = n10379 ^ n4606;
  assign n10381 = n10015 & ~n10229;
  assign n10382 = n10381 ^ n10017;
  assign n10383 = n10382 ^ n10379;
  assign n10384 = n10380 & n10383;
  assign n10385 = n10384 ^ n4606;
  assign n10386 = n10385 ^ n4362;
  assign n10387 = n10021 & ~n10229;
  assign n10388 = n10387 ^ n10024;
  assign n10389 = n10388 ^ n10385;
  assign n10390 = n10386 & ~n10389;
  assign n10391 = n10390 ^ n4362;
  assign n10392 = n10391 ^ n4133;
  assign n10393 = n10028 & ~n10229;
  assign n10394 = n10393 ^ n10031;
  assign n10395 = n10394 ^ n10391;
  assign n10396 = n10392 & n10395;
  assign n10397 = n10396 ^ n4133;
  assign n10398 = n10397 ^ n3882;
  assign n10399 = n10035 & ~n10229;
  assign n10400 = n10399 ^ n10037;
  assign n10401 = n10400 ^ n10397;
  assign n10402 = n10398 & ~n10401;
  assign n10403 = n10402 ^ n3882;
  assign n10404 = n10403 ^ n3634;
  assign n10405 = n10040 ^ n3882;
  assign n10406 = ~n10229 & n10405;
  assign n10407 = n10406 ^ n9881;
  assign n10408 = n10407 ^ n10403;
  assign n10409 = ~n10404 & n10408;
  assign n10410 = n10409 ^ n3634;
  assign n10411 = n10410 ^ n3397;
  assign n10412 = n10043 ^ n3634;
  assign n10413 = ~n10229 & ~n10412;
  assign n10414 = n10413 ^ n9878;
  assign n10415 = n10414 ^ n10410;
  assign n10416 = ~n10411 & n10415;
  assign n10417 = n10416 ^ n3397;
  assign n10418 = n10417 ^ n3177;
  assign n10419 = ~n10047 & ~n10229;
  assign n10420 = n10419 ^ n10049;
  assign n10421 = n10420 ^ n10417;
  assign n10422 = n10418 & n10421;
  assign n10423 = n10422 ^ n3177;
  assign n10424 = n10423 ^ n2980;
  assign n10425 = n10053 & ~n10229;
  assign n10426 = n10425 ^ n10056;
  assign n10427 = n10426 ^ n10423;
  assign n10428 = n10424 & ~n10427;
  assign n10429 = n10428 ^ n2980;
  assign n10430 = n10429 ^ n2782;
  assign n10431 = n10060 & ~n10229;
  assign n10432 = n10431 ^ n10063;
  assign n10433 = n10432 ^ n10429;
  assign n10434 = n10430 & n10433;
  assign n10435 = n10434 ^ n2782;
  assign n10436 = n10435 ^ n10248;
  assign n10437 = n10249 & ~n10436;
  assign n10438 = n10437 ^ n2583;
  assign n10439 = n10438 ^ n10245;
  assign n10440 = ~n10246 & n10439;
  assign n10441 = n10440 ^ n2374;
  assign n10442 = n10441 ^ n2194;
  assign n10443 = n10079 & ~n10229;
  assign n10444 = n10443 ^ n10081;
  assign n10445 = n10444 ^ n10441;
  assign n10446 = ~n10442 & ~n10445;
  assign n10447 = n10446 ^ n2194;
  assign n10448 = n10447 ^ n2011;
  assign n10449 = ~n10085 & ~n10229;
  assign n10450 = n10449 ^ n10087;
  assign n10451 = n10450 ^ n10447;
  assign n10452 = ~n10448 & ~n10451;
  assign n10453 = n10452 ^ n2011;
  assign n10454 = n10453 ^ n1804;
  assign n10455 = ~n10091 & ~n10229;
  assign n10456 = n10455 ^ n10093;
  assign n10457 = n10456 ^ n10453;
  assign n10458 = n10454 & ~n10457;
  assign n10459 = n10458 ^ n1804;
  assign n10460 = n10459 ^ n1621;
  assign n10461 = n10097 & ~n10229;
  assign n10462 = n10461 ^ n10099;
  assign n10463 = n10462 ^ n10459;
  assign n10464 = n10460 & n10463;
  assign n10465 = n10464 ^ n1621;
  assign n10466 = n10465 ^ n10242;
  assign n10467 = n10243 & ~n10466;
  assign n10468 = n10467 ^ n1458;
  assign n10469 = n10468 ^ n10239;
  assign n10470 = ~n10240 & n10469;
  assign n10471 = n10470 ^ n1299;
  assign n10472 = n10471 ^ n10236;
  assign n10473 = n10237 & ~n10472;
  assign n10474 = n10473 ^ n1158;
  assign n10475 = n10474 ^ n10232;
  assign n10476 = ~n10233 & n10475;
  assign n10477 = n10476 ^ n1027;
  assign n10478 = n10477 ^ n905;
  assign n10479 = n10121 & ~n10229;
  assign n10480 = n10479 ^ n10123;
  assign n10481 = n10480 ^ n10477;
  assign n10482 = n10478 & ~n10481;
  assign n10483 = n10482 ^ n905;
  assign n10484 = n10483 ^ n803;
  assign n10485 = n10127 & ~n10229;
  assign n10486 = n10485 ^ n10129;
  assign n10487 = n10486 ^ n10483;
  assign n10488 = n10484 & n10487;
  assign n10489 = n10488 ^ n803;
  assign n10490 = n10489 ^ n707;
  assign n10491 = n10133 & ~n10229;
  assign n10492 = n10491 ^ n10135;
  assign n10493 = n10492 ^ n10489;
  assign n10494 = ~n10490 & ~n10493;
  assign n10495 = n10494 ^ n707;
  assign n10496 = n10495 ^ n608;
  assign n10497 = ~n10139 & ~n10229;
  assign n10498 = n10497 ^ n10141;
  assign n10499 = n10498 ^ n10495;
  assign n10500 = ~n10496 & ~n10499;
  assign n10501 = n10500 ^ n608;
  assign n10502 = n10501 ^ n514;
  assign n10503 = ~n10145 & ~n10229;
  assign n10504 = n10503 ^ n10147;
  assign n10505 = n10504 ^ n10501;
  assign n10506 = n10502 & ~n10505;
  assign n10507 = n10506 ^ n514;
  assign n10508 = n10507 ^ n436;
  assign n10509 = n10151 & ~n10229;
  assign n10510 = n10509 ^ n10154;
  assign n10511 = n10510 ^ n10507;
  assign n10512 = n10508 & n10511;
  assign n10513 = n10512 ^ n436;
  assign n10514 = n10513 ^ n363;
  assign n10515 = n10158 & ~n10229;
  assign n10516 = n10515 ^ n10161;
  assign n10517 = n10516 ^ n10513;
  assign n10518 = n10514 & ~n10517;
  assign n10519 = n10518 ^ n363;
  assign n10520 = n10519 ^ n300;
  assign n10521 = n132 & n10197;
  assign n10522 = ~n10228 & ~n10521;
  assign n10523 = ~n133 & ~n10522;
  assign n10524 = n133 & ~n10199;
  assign n10525 = n10198 & n10524;
  assign n10526 = n129 & ~n10227;
  assign n10527 = ~n1287 & ~n10526;
  assign n10528 = n9869 & ~n10527;
  assign n10529 = n10197 & n10528;
  assign n10530 = ~n10203 & ~n10529;
  assign n10531 = ~n10525 & n10530;
  assign n10532 = ~n10523 & n10531;
  assign n10533 = ~n133 & ~n10200;
  assign n10534 = n10203 & ~n10533;
  assign n10535 = ~n10532 & ~n10534;
  assign n10536 = n10228 ^ n10203;
  assign n10537 = n133 & ~n10536;
  assign n10538 = n10537 ^ n10203;
  assign n10539 = n10538 ^ n10197;
  assign n10540 = n10538 ^ n132;
  assign n10541 = n10540 ^ n132;
  assign n10542 = n1292 & n10203;
  assign n10543 = n10542 ^ n132;
  assign n10544 = n10541 & ~n10543;
  assign n10545 = n10544 ^ n132;
  assign n10546 = ~n10539 & n10545;
  assign n10547 = n10546 ^ n10197;
  assign n10548 = ~n9869 & n10547;
  assign n10549 = ~n10535 & ~n10548;
  assign n10550 = n10197 ^ n132;
  assign n10551 = ~n10229 & n10550;
  assign n10552 = n10551 ^ n9869;
  assign n10553 = ~n10549 & ~n10552;
  assign n10554 = ~n133 & n10553;
  assign n10557 = n10165 & ~n10229;
  assign n10558 = n10557 ^ n10167;
  assign n10559 = n10558 ^ n10519;
  assign n10560 = n10520 & ~n10559;
  assign n10561 = n10560 ^ n300;
  assign n10562 = n10561 ^ n243;
  assign n10563 = n10171 & ~n10229;
  assign n10564 = n10563 ^ n10174;
  assign n10565 = n10564 ^ n10561;
  assign n10566 = n10562 & ~n10565;
  assign n10567 = n10566 ^ n243;
  assign n10568 = n10567 ^ n210;
  assign n10569 = n10178 & ~n10229;
  assign n10570 = n10569 ^ n10181;
  assign n10571 = n10570 ^ n10567;
  assign n10572 = n10568 & n10571;
  assign n10573 = n10572 ^ n210;
  assign n10574 = n10573 ^ n147;
  assign n10575 = n10185 & ~n10229;
  assign n10576 = n10575 ^ n10188;
  assign n10577 = n10576 ^ n10573;
  assign n10578 = ~n10574 & ~n10577;
  assign n10579 = n10578 ^ n147;
  assign n10555 = ~n10192 & ~n10229;
  assign n10556 = n10555 ^ n10194;
  assign n10580 = n10579 ^ n10556;
  assign n10581 = n10556 ^ n132;
  assign n10582 = n10580 & n10581;
  assign n10583 = n10582 ^ n10556;
  assign n10584 = ~n10549 & n10583;
  assign n10585 = ~n10554 & ~n10584;
  assign n10586 = n10520 & n10585;
  assign n10587 = n10586 ^ n10558;
  assign n10588 = n10587 ^ n243;
  assign n10589 = n10514 & n10585;
  assign n10590 = n10589 ^ n10516;
  assign n10591 = n10590 ^ n300;
  assign n10592 = n10468 ^ n1299;
  assign n10593 = n10585 & n10592;
  assign n10594 = n10593 ^ n10239;
  assign n10595 = n10594 ^ n1158;
  assign n10596 = n10465 ^ n1458;
  assign n10597 = n10585 & n10596;
  assign n10598 = n10597 ^ n10242;
  assign n10599 = n10598 ^ n1299;
  assign n10600 = ~n10404 & n10585;
  assign n10601 = n10600 ^ n10407;
  assign n10602 = n10601 ^ n3397;
  assign n10603 = n10398 & n10585;
  assign n10604 = n10603 ^ n10400;
  assign n10605 = n10604 ^ n3634;
  assign n10606 = n10374 & n10585;
  assign n10607 = n10606 ^ n10376;
  assign n10608 = n10607 ^ n4606;
  assign n10609 = n10368 & n10585;
  assign n10610 = n10609 ^ n10370;
  assign n10611 = n10610 ^ n4851;
  assign n10612 = n10350 & n10585;
  assign n10613 = n10612 ^ n10352;
  assign n10614 = n10613 ^ n5625;
  assign n10615 = n10344 & n10585;
  assign n10616 = n10615 ^ n10346;
  assign n10617 = n10616 ^ n5905;
  assign n10618 = n10585 ^ x26;
  assign n10619 = n10618 ^ x26;
  assign n10620 = ~x24 & ~x25;
  assign n10621 = n10229 & n10620;
  assign n10622 = ~x26 & n10621;
  assign n10623 = n10622 ^ n10229;
  assign n10624 = n10623 ^ x26;
  assign n10625 = ~n10619 & ~n10624;
  assign n10626 = n10625 ^ x26;
  assign n10627 = ~x27 & n10626;
  assign n10628 = n10620 ^ x26;
  assign n10629 = ~x26 & ~n10628;
  assign n10630 = n10629 ^ n10229;
  assign n10631 = n10630 ^ x26;
  assign n10632 = x27 & n10585;
  assign n10633 = n10632 ^ n10229;
  assign n10634 = n10631 & ~n10633;
  assign n10635 = n10634 ^ n10229;
  assign n10636 = ~n10627 & n10635;
  assign n10637 = n10636 ^ n9867;
  assign n10638 = n10251 ^ n10229;
  assign n10639 = n10585 & ~n10638;
  assign n10640 = n10639 ^ n10229;
  assign n10641 = n10640 ^ x28;
  assign n10642 = n10641 ^ n10636;
  assign n10643 = n10637 & n10642;
  assign n10644 = n10643 ^ n9867;
  assign n10645 = n10644 ^ n9502;
  assign n10647 = ~x28 & n10251;
  assign n10648 = n10647 ^ n9867;
  assign n10649 = n10648 ^ n10250;
  assign n10650 = n10229 & ~n10649;
  assign n10651 = n10650 ^ n10250;
  assign n10646 = ~x28 & ~n10229;
  assign n10652 = n10651 ^ n10646;
  assign n10653 = n10251 ^ n9867;
  assign n10654 = n10653 ^ n10651;
  assign n10655 = n10651 ^ n10585;
  assign n10656 = ~n10651 & ~n10655;
  assign n10657 = n10656 ^ n10651;
  assign n10658 = ~n10654 & ~n10657;
  assign n10659 = n10658 ^ n10656;
  assign n10660 = n10659 ^ n10651;
  assign n10661 = n10660 ^ n10585;
  assign n10662 = n10652 & ~n10661;
  assign n10663 = n10662 ^ n10646;
  assign n10664 = n10663 ^ x29;
  assign n10665 = n10664 ^ n10644;
  assign n10666 = n10645 & ~n10665;
  assign n10667 = n10666 ^ n9502;
  assign n10668 = n10667 ^ n9129;
  assign n10669 = n10262 & n10585;
  assign n10670 = n10669 ^ n10266;
  assign n10671 = n10670 ^ n10667;
  assign n10672 = n10668 & n10671;
  assign n10673 = n10672 ^ n9129;
  assign n10674 = n10673 ^ n8769;
  assign n10675 = n10270 & n10585;
  assign n10676 = n10675 ^ n10292;
  assign n10677 = n10676 ^ n10673;
  assign n10678 = n10674 & ~n10677;
  assign n10679 = n10678 ^ n8769;
  assign n10680 = n10679 ^ n8422;
  assign n10681 = n10296 & n10585;
  assign n10682 = n10681 ^ n10298;
  assign n10683 = n10682 ^ n10679;
  assign n10684 = n10680 & n10683;
  assign n10685 = n10684 ^ n8422;
  assign n10686 = n10685 ^ n8083;
  assign n10687 = n10302 & n10585;
  assign n10688 = n10687 ^ n10304;
  assign n10689 = n10688 ^ n10685;
  assign n10690 = n10686 & ~n10689;
  assign n10691 = n10690 ^ n8083;
  assign n10692 = n10691 ^ n7777;
  assign n10693 = n10308 & n10585;
  assign n10694 = n10693 ^ n10310;
  assign n10695 = n10694 ^ n10691;
  assign n10696 = n10692 & n10695;
  assign n10697 = n10696 ^ n7777;
  assign n10698 = n10697 ^ n7463;
  assign n10699 = n10314 & n10585;
  assign n10700 = n10699 ^ n10316;
  assign n10701 = n10700 ^ n10697;
  assign n10702 = n10698 & ~n10701;
  assign n10703 = n10702 ^ n7463;
  assign n10704 = n10703 ^ n7135;
  assign n10705 = n10320 & n10585;
  assign n10706 = n10705 ^ n10322;
  assign n10707 = n10706 ^ n10703;
  assign n10708 = n10704 & n10707;
  assign n10709 = n10708 ^ n7135;
  assign n10710 = n10709 ^ n6802;
  assign n10711 = n10326 & n10585;
  assign n10712 = n10711 ^ n10328;
  assign n10713 = n10712 ^ n10709;
  assign n10714 = n10710 & ~n10713;
  assign n10715 = n10714 ^ n6802;
  assign n10716 = n10715 ^ n6479;
  assign n10717 = n10332 & n10585;
  assign n10718 = n10717 ^ n10334;
  assign n10719 = n10718 ^ n10715;
  assign n10720 = n10716 & n10719;
  assign n10721 = n10720 ^ n6479;
  assign n10722 = n10721 ^ n6181;
  assign n10723 = n10338 & n10585;
  assign n10724 = n10723 ^ n10340;
  assign n10725 = n10724 ^ n10721;
  assign n10726 = n10722 & ~n10725;
  assign n10727 = n10726 ^ n6181;
  assign n10728 = n10727 ^ n10616;
  assign n10729 = ~n10617 & n10728;
  assign n10730 = n10729 ^ n5905;
  assign n10731 = n10730 ^ n10613;
  assign n10732 = n10614 & ~n10731;
  assign n10733 = n10732 ^ n5625;
  assign n10734 = n10733 ^ n5363;
  assign n10735 = n10356 & n10585;
  assign n10736 = n10735 ^ n10358;
  assign n10737 = n10736 ^ n10733;
  assign n10738 = n10734 & ~n10737;
  assign n10739 = n10738 ^ n5363;
  assign n10740 = n10739 ^ n5108;
  assign n10741 = n10362 & n10585;
  assign n10742 = n10741 ^ n10364;
  assign n10743 = n10742 ^ n10739;
  assign n10744 = n10740 & ~n10743;
  assign n10745 = n10744 ^ n5108;
  assign n10746 = n10745 ^ n10610;
  assign n10747 = ~n10611 & n10746;
  assign n10748 = n10747 ^ n4851;
  assign n10749 = n10748 ^ n10607;
  assign n10750 = n10608 & ~n10749;
  assign n10751 = n10750 ^ n4606;
  assign n10752 = n10751 ^ n4362;
  assign n10753 = n10380 & n10585;
  assign n10754 = n10753 ^ n10382;
  assign n10755 = n10754 ^ n10751;
  assign n10756 = n10752 & n10755;
  assign n10757 = n10756 ^ n4362;
  assign n10758 = n10757 ^ n4133;
  assign n10759 = n10386 & n10585;
  assign n10760 = n10759 ^ n10388;
  assign n10761 = n10760 ^ n10757;
  assign n10762 = n10758 & ~n10761;
  assign n10763 = n10762 ^ n4133;
  assign n10764 = n10763 ^ n3882;
  assign n10765 = n10392 & n10585;
  assign n10766 = n10765 ^ n10394;
  assign n10767 = n10766 ^ n10763;
  assign n10768 = n10764 & n10767;
  assign n10769 = n10768 ^ n3882;
  assign n10770 = n10769 ^ n10604;
  assign n10771 = ~n10605 & ~n10770;
  assign n10772 = n10771 ^ n3634;
  assign n10773 = n10772 ^ n10601;
  assign n10774 = ~n10602 & ~n10773;
  assign n10775 = n10774 ^ n3397;
  assign n10776 = n10775 ^ n3177;
  assign n10777 = ~n10411 & n10585;
  assign n10778 = n10777 ^ n10414;
  assign n10779 = n10778 ^ n10775;
  assign n10780 = n10776 & ~n10779;
  assign n10781 = n10780 ^ n3177;
  assign n10782 = n10781 ^ n2980;
  assign n10783 = n10418 & n10585;
  assign n10784 = n10783 ^ n10420;
  assign n10785 = n10784 ^ n10781;
  assign n10786 = n10782 & n10785;
  assign n10787 = n10786 ^ n2980;
  assign n10788 = n10787 ^ n2782;
  assign n10789 = n10424 & n10585;
  assign n10790 = n10789 ^ n10426;
  assign n10791 = n10790 ^ n10787;
  assign n10792 = n10788 & ~n10791;
  assign n10793 = n10792 ^ n2782;
  assign n10794 = n10793 ^ n2583;
  assign n10795 = n10430 & n10585;
  assign n10796 = n10795 ^ n10432;
  assign n10797 = n10796 ^ n10793;
  assign n10798 = n10794 & n10797;
  assign n10799 = n10798 ^ n2583;
  assign n10800 = n10799 ^ n2374;
  assign n10801 = n10435 ^ n2583;
  assign n10802 = n10585 & n10801;
  assign n10803 = n10802 ^ n10248;
  assign n10804 = n10803 ^ n10799;
  assign n10805 = n10800 & ~n10804;
  assign n10806 = n10805 ^ n2374;
  assign n10807 = n10806 ^ n2194;
  assign n10808 = n10438 ^ n2374;
  assign n10809 = n10585 & n10808;
  assign n10810 = n10809 ^ n10245;
  assign n10811 = n10810 ^ n10806;
  assign n10812 = ~n10807 & n10811;
  assign n10813 = n10812 ^ n2194;
  assign n10814 = n10813 ^ n2011;
  assign n10815 = ~n10442 & n10585;
  assign n10816 = n10815 ^ n10444;
  assign n10817 = n10816 ^ n10813;
  assign n10818 = ~n10814 & n10817;
  assign n10819 = n10818 ^ n2011;
  assign n10820 = n10819 ^ n1804;
  assign n10821 = ~n10448 & n10585;
  assign n10822 = n10821 ^ n10450;
  assign n10823 = n10822 ^ n10819;
  assign n10824 = n10820 & n10823;
  assign n10825 = n10824 ^ n1804;
  assign n10826 = n10825 ^ n1621;
  assign n10827 = n10454 & n10585;
  assign n10828 = n10827 ^ n10456;
  assign n10829 = n10828 ^ n10825;
  assign n10830 = n10826 & ~n10829;
  assign n10831 = n10830 ^ n1621;
  assign n10832 = n10831 ^ n1458;
  assign n10833 = n10460 & n10585;
  assign n10834 = n10833 ^ n10462;
  assign n10835 = n10834 ^ n10831;
  assign n10836 = n10832 & n10835;
  assign n10837 = n10836 ^ n1458;
  assign n10838 = n10837 ^ n10598;
  assign n10839 = n10599 & ~n10838;
  assign n10840 = n10839 ^ n1299;
  assign n10841 = n10840 ^ n10594;
  assign n10842 = ~n10595 & n10841;
  assign n10843 = n10842 ^ n1158;
  assign n10844 = n10843 ^ n1027;
  assign n10845 = n10471 ^ n1158;
  assign n10846 = n10585 & n10845;
  assign n10847 = n10846 ^ n10236;
  assign n10848 = n10847 ^ n10843;
  assign n10849 = n10844 & ~n10848;
  assign n10850 = n10849 ^ n1027;
  assign n10851 = n10850 ^ n905;
  assign n10852 = n10474 ^ n1027;
  assign n10853 = n10585 & n10852;
  assign n10854 = n10853 ^ n10232;
  assign n10855 = n10854 ^ n10850;
  assign n10856 = n10851 & n10855;
  assign n10857 = n10856 ^ n905;
  assign n10858 = n10857 ^ n803;
  assign n10859 = n10478 & n10585;
  assign n10860 = n10859 ^ n10480;
  assign n10861 = n10860 ^ n10857;
  assign n10862 = n10858 & ~n10861;
  assign n10863 = n10862 ^ n803;
  assign n10864 = n10863 ^ n707;
  assign n10865 = n10484 & n10585;
  assign n10866 = n10865 ^ n10486;
  assign n10867 = n10866 ^ n10863;
  assign n10868 = ~n10864 & n10867;
  assign n10869 = n10868 ^ n707;
  assign n10870 = n10869 ^ n608;
  assign n10871 = ~n10490 & n10585;
  assign n10872 = n10871 ^ n10492;
  assign n10873 = n10872 ^ n10869;
  assign n10874 = ~n10870 & n10873;
  assign n10875 = n10874 ^ n608;
  assign n10876 = n10875 ^ n514;
  assign n10877 = ~n10496 & n10585;
  assign n10878 = n10877 ^ n10498;
  assign n10879 = n10878 ^ n10875;
  assign n10880 = n10876 & n10879;
  assign n10881 = n10880 ^ n514;
  assign n10882 = n10881 ^ n436;
  assign n10883 = n10502 & n10585;
  assign n10884 = n10883 ^ n10504;
  assign n10885 = n10884 ^ n10881;
  assign n10886 = n10882 & ~n10885;
  assign n10887 = n10886 ^ n436;
  assign n10888 = n10887 ^ n363;
  assign n10889 = n10508 & n10585;
  assign n10890 = n10889 ^ n10510;
  assign n10891 = n10890 ^ n10887;
  assign n10892 = n10888 & n10891;
  assign n10893 = n10892 ^ n363;
  assign n10894 = n10893 ^ n10590;
  assign n10895 = n10591 & ~n10894;
  assign n10896 = n10895 ^ n300;
  assign n10897 = n10896 ^ n10587;
  assign n10898 = n10588 & ~n10897;
  assign n10899 = n10898 ^ n243;
  assign n10900 = n10899 ^ n210;
  assign n10901 = n10562 & n10585;
  assign n10902 = n10901 ^ n10564;
  assign n10903 = n10902 ^ n10899;
  assign n10904 = n10900 & ~n10903;
  assign n10905 = n10904 ^ n210;
  assign n10906 = n10905 ^ n147;
  assign n10907 = n10579 ^ n132;
  assign n10908 = n10585 & n10907;
  assign n10909 = n10908 ^ n10556;
  assign n10910 = ~n133 & n10909;
  assign n10911 = n10568 & n10585;
  assign n10912 = n10911 ^ n10570;
  assign n10913 = n10912 ^ n10905;
  assign n10914 = ~n10906 & n10913;
  assign n10915 = n10914 ^ n147;
  assign n10916 = n10915 ^ n132;
  assign n10917 = ~n10574 & n10585;
  assign n10918 = n10917 ^ n10576;
  assign n10919 = n10918 ^ n10915;
  assign n10920 = n10916 & n10919;
  assign n10921 = n10920 ^ n132;
  assign n10922 = ~n10910 & ~n10921;
  assign n10923 = n132 & n10579;
  assign n10924 = n10549 & ~n10552;
  assign n10925 = ~n10556 & ~n10924;
  assign n10926 = ~n10923 & n10925;
  assign n10927 = n10552 ^ n132;
  assign n10928 = n10927 ^ n10579;
  assign n10929 = n10928 ^ n10552;
  assign n10930 = n10579 ^ n10552;
  assign n10931 = n10930 ^ n10579;
  assign n10932 = n10580 ^ n10579;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = n10933 ^ n10579;
  assign n10935 = n10929 & n10934;
  assign n10936 = n10935 ^ n10927;
  assign n10937 = ~n10926 & ~n10936;
  assign n10938 = ~n133 & ~n10937;
  assign n10939 = n10556 & n10579;
  assign n10940 = ~n10552 & ~n10939;
  assign n10941 = ~n132 & ~n10940;
  assign n10942 = n10549 & n10556;
  assign n10943 = n10923 & ~n10942;
  assign n10944 = ~n132 & ~n10556;
  assign n10945 = ~n10552 & ~n10944;
  assign n10946 = ~n10579 & ~n10945;
  assign n10947 = n132 & n10556;
  assign n10948 = ~n10552 & n10947;
  assign n10949 = n133 & ~n10948;
  assign n10950 = ~n10946 & n10949;
  assign n10951 = ~n10943 & n10950;
  assign n10952 = ~n10941 & n10951;
  assign n10953 = n10553 & n10556;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = ~n10938 & n10954;
  assign n10956 = ~n10922 & ~n10955;
  assign n10957 = ~n10906 & ~n10956;
  assign n10958 = n10957 ^ n10912;
  assign n10959 = ~n132 & ~n10958;
  assign n10960 = n10882 & ~n10956;
  assign n10961 = n10960 ^ n10884;
  assign n10962 = n363 & n10961;
  assign n10963 = n10840 ^ n1158;
  assign n10964 = ~n10956 & n10963;
  assign n10965 = n10964 ^ n10594;
  assign n10966 = n10965 ^ n1027;
  assign n10967 = n10837 ^ n1299;
  assign n10968 = ~n10956 & n10967;
  assign n10969 = n10968 ^ n10598;
  assign n10970 = n10969 ^ n1158;
  assign n10971 = n10740 & ~n10956;
  assign n10972 = n10971 ^ n10742;
  assign n10973 = n10972 ^ n4851;
  assign n10974 = n10730 ^ n5625;
  assign n10975 = ~n10956 & n10974;
  assign n10976 = n10975 ^ n10613;
  assign n10977 = ~n5363 & ~n10976;
  assign n10978 = n10727 ^ n5905;
  assign n10979 = ~n10956 & n10978;
  assign n10980 = n10979 ^ n10616;
  assign n10981 = ~n5625 & n10980;
  assign n10982 = ~n10977 & ~n10981;
  assign n10983 = n10698 & ~n10956;
  assign n10984 = n10983 ^ n10700;
  assign n10985 = n10984 ^ n7135;
  assign n10986 = n10692 & ~n10956;
  assign n10987 = n10986 ^ n10694;
  assign n10988 = n10987 ^ n7463;
  assign n10989 = n10686 & ~n10956;
  assign n10990 = n10989 ^ n10688;
  assign n10991 = n10990 ^ n7777;
  assign n10992 = n10680 & ~n10956;
  assign n10993 = n10992 ^ n10682;
  assign n10994 = n10993 ^ n8083;
  assign n10995 = n10637 & ~n10956;
  assign n10996 = n10995 ^ n10641;
  assign n10997 = n10996 ^ n9502;
  assign n11020 = x26 & n10585;
  assign n11021 = ~x22 & ~x23;
  assign n11022 = ~x24 & n11021;
  assign n11023 = n10585 & n11022;
  assign n11024 = ~n11020 & ~n11023;
  assign n11025 = n10620 & ~n10956;
  assign n11026 = ~x26 & ~n11025;
  assign n11027 = x25 & n10585;
  assign n11028 = ~n10955 & n11027;
  assign n11029 = n11028 ^ n11025;
  assign n11030 = n11026 ^ n10922;
  assign n11031 = ~n11029 & n11030;
  assign n11032 = n11031 ^ n10922;
  assign n11033 = n11026 & n11032;
  assign n11034 = n11024 & ~n11033;
  assign n11036 = x26 ^ x25;
  assign n11037 = n11036 ^ n11022;
  assign n11038 = n11037 ^ x26;
  assign n11035 = n10956 ^ x26;
  assign n11039 = n11038 ^ n11035;
  assign n11040 = n11022 ^ n10956;
  assign n11041 = n11040 ^ x26;
  assign n11042 = n11041 ^ x26;
  assign n11043 = ~n11037 & ~n11042;
  assign n11044 = n11043 ^ n11037;
  assign n11045 = n11041 & ~n11044;
  assign n11046 = n11045 ^ x26;
  assign n11047 = n11039 & ~n11046;
  assign n11048 = n11047 ^ n11043;
  assign n11049 = n11048 ^ x26;
  assign n11050 = n11049 ^ n11035;
  assign n11051 = n11034 & n11050;
  assign n11052 = ~n10229 & ~n11051;
  assign n11053 = n10956 ^ x25;
  assign n11054 = ~n11040 & ~n11053;
  assign n11055 = n11054 ^ x25;
  assign n11056 = n11020 & ~n11055;
  assign n11057 = n10956 ^ n10620;
  assign n11058 = n11057 ^ x26;
  assign n11061 = ~n10585 & n11021;
  assign n11059 = ~n10585 & ~n11022;
  assign n11060 = x25 & n11059;
  assign n11062 = n11061 ^ n11060;
  assign n11063 = n11060 ^ n10956;
  assign n11064 = n11063 ^ n11060;
  assign n11065 = ~n11062 & n11064;
  assign n11066 = n11065 ^ n11060;
  assign n11067 = n11066 ^ n11057;
  assign n11068 = n11058 & n11067;
  assign n11069 = n11068 ^ n11065;
  assign n11070 = n11069 ^ n11060;
  assign n11071 = n11070 ^ x26;
  assign n11072 = ~n11057 & n11071;
  assign n11073 = n11072 ^ n11057;
  assign n11074 = ~n11056 & n11073;
  assign n11075 = ~n11052 & n11074;
  assign n10999 = n10585 ^ n10229;
  assign n11000 = n10999 ^ n10585;
  assign n11001 = n11000 ^ n10999;
  assign n11002 = n10999 ^ n10620;
  assign n11003 = ~n11001 & ~n11002;
  assign n11004 = n11003 ^ n10999;
  assign n11005 = ~x26 & ~n11004;
  assign n11006 = n11005 ^ n10999;
  assign n10998 = ~x26 & n10585;
  assign n11007 = n11006 ^ n10998;
  assign n11008 = n10620 ^ n10229;
  assign n11009 = n11008 ^ n11006;
  assign n11010 = n11006 ^ n10956;
  assign n11011 = n11006 & ~n11010;
  assign n11012 = n11011 ^ n11006;
  assign n11013 = n11009 & n11012;
  assign n11014 = n11013 ^ n11011;
  assign n11015 = n11014 ^ n11006;
  assign n11016 = n11015 ^ n10956;
  assign n11017 = ~n11007 & ~n11016;
  assign n11018 = n11017 ^ n10998;
  assign n11019 = n11018 ^ x27;
  assign n11076 = n11075 ^ n11019;
  assign n11077 = n11075 ^ n9867;
  assign n11078 = ~n11076 & n11077;
  assign n11079 = n11078 ^ n9867;
  assign n11080 = n11079 ^ n10996;
  assign n11081 = ~n10997 & n11080;
  assign n11082 = n11081 ^ n9502;
  assign n11083 = n11082 ^ n9129;
  assign n11084 = n10645 & ~n10956;
  assign n11085 = n11084 ^ n10664;
  assign n11086 = n11085 ^ n11082;
  assign n11087 = n11083 & ~n11086;
  assign n11088 = n11087 ^ n9129;
  assign n11089 = n11088 ^ n8769;
  assign n11090 = n10668 & ~n10956;
  assign n11091 = n11090 ^ n10670;
  assign n11092 = n11091 ^ n11088;
  assign n11093 = n11089 & n11092;
  assign n11094 = n11093 ^ n8769;
  assign n11095 = n11094 ^ n8422;
  assign n11096 = n10674 & ~n10956;
  assign n11097 = n11096 ^ n10676;
  assign n11098 = n11097 ^ n11094;
  assign n11099 = n11095 & ~n11098;
  assign n11100 = n11099 ^ n8422;
  assign n11101 = n11100 ^ n10993;
  assign n11102 = ~n10994 & n11101;
  assign n11103 = n11102 ^ n8083;
  assign n11104 = n11103 ^ n10990;
  assign n11105 = n10991 & ~n11104;
  assign n11106 = n11105 ^ n7777;
  assign n11107 = n11106 ^ n10987;
  assign n11108 = ~n10988 & n11107;
  assign n11109 = n11108 ^ n7463;
  assign n11110 = n11109 ^ n10984;
  assign n11111 = n10985 & ~n11110;
  assign n11112 = n11111 ^ n7135;
  assign n11113 = n11112 ^ n6802;
  assign n11114 = n10704 & ~n10956;
  assign n11115 = n11114 ^ n10706;
  assign n11116 = n11115 ^ n11112;
  assign n11117 = n11113 & n11116;
  assign n11118 = n11117 ^ n6802;
  assign n11119 = n11118 ^ n6479;
  assign n11120 = n10710 & ~n10956;
  assign n11121 = n11120 ^ n10712;
  assign n11122 = n11121 ^ n11118;
  assign n11123 = n11119 & ~n11122;
  assign n11124 = n11123 ^ n6479;
  assign n11125 = n11124 ^ n6181;
  assign n11126 = n10716 & ~n10956;
  assign n11127 = n11126 ^ n10718;
  assign n11128 = n11127 ^ n11124;
  assign n11129 = n11125 & n11128;
  assign n11130 = n11129 ^ n6181;
  assign n11131 = n11130 ^ n5905;
  assign n11132 = n10722 & ~n10956;
  assign n11133 = n11132 ^ n10724;
  assign n11134 = n11133 ^ n11130;
  assign n11135 = n11131 & ~n11134;
  assign n11136 = n11135 ^ n5905;
  assign n11137 = n10982 & n11136;
  assign n11138 = n5625 & ~n10980;
  assign n11139 = ~n10977 & n11138;
  assign n11140 = n5363 & n10976;
  assign n11141 = n10734 & ~n10956;
  assign n11142 = n11141 ^ n10736;
  assign n11143 = n5108 & n11142;
  assign n11144 = ~n11140 & ~n11143;
  assign n11145 = ~n11139 & n11144;
  assign n11146 = ~n11137 & n11145;
  assign n11147 = n11146 ^ n10972;
  assign n11148 = n11147 ^ n10972;
  assign n11149 = ~n5108 & ~n11142;
  assign n11150 = n11149 ^ n10972;
  assign n11151 = n11150 ^ n10972;
  assign n11152 = ~n11148 & ~n11151;
  assign n11153 = n11152 ^ n10972;
  assign n11154 = n10973 & ~n11153;
  assign n11155 = n11154 ^ n4851;
  assign n11156 = n4606 & n11155;
  assign n11157 = n10748 ^ n4606;
  assign n11158 = ~n10956 & n11157;
  assign n11159 = n11158 ^ n10607;
  assign n11160 = n11156 & n11159;
  assign n11161 = n10745 ^ n4851;
  assign n11162 = ~n10956 & n11161;
  assign n11163 = n11162 ^ n10610;
  assign n11164 = n11163 ^ n4362;
  assign n11165 = n11159 ^ n4606;
  assign n11166 = n11163 ^ n4606;
  assign n11167 = n11166 ^ n4606;
  assign n11168 = ~n11165 & ~n11167;
  assign n11169 = n11168 ^ n4606;
  assign n11170 = ~n11164 & ~n11169;
  assign n11171 = n11170 ^ n4362;
  assign n11172 = n11155 & n11171;
  assign n11173 = n11159 ^ n4362;
  assign n11174 = n11163 ^ n11159;
  assign n11175 = n11174 ^ n11159;
  assign n11176 = n11165 ^ n11159;
  assign n11177 = ~n11175 & n11176;
  assign n11178 = n11177 ^ n11159;
  assign n11179 = n11173 & ~n11178;
  assign n11180 = n11179 ^ n4362;
  assign n11181 = ~n11172 & ~n11180;
  assign n11182 = ~n11160 & n11181;
  assign n11183 = n10752 & ~n10956;
  assign n11184 = n11183 ^ n10754;
  assign n11185 = ~n4133 & n11184;
  assign n11186 = n10758 & ~n10956;
  assign n11187 = n11186 ^ n10760;
  assign n11188 = ~n3882 & ~n11187;
  assign n11189 = ~n11185 & ~n11188;
  assign n11190 = ~n11182 & n11189;
  assign n11191 = n11187 ^ n3882;
  assign n11192 = n4133 & ~n11184;
  assign n11193 = n11192 ^ n11187;
  assign n11194 = n11191 & ~n11193;
  assign n11195 = n11194 ^ n3882;
  assign n11196 = ~n11190 & ~n11195;
  assign n11197 = n11196 ^ n3634;
  assign n11198 = n10764 & ~n10956;
  assign n11199 = n11198 ^ n10766;
  assign n11200 = n11199 ^ n11196;
  assign n11201 = n11197 & ~n11200;
  assign n11202 = n11201 ^ n3634;
  assign n11203 = n11202 ^ n3397;
  assign n11204 = n10769 ^ n3634;
  assign n11205 = ~n10956 & ~n11204;
  assign n11206 = n11205 ^ n10604;
  assign n11207 = n11206 ^ n11202;
  assign n11208 = ~n11203 & n11207;
  assign n11209 = n11208 ^ n3397;
  assign n11210 = n11209 ^ n3177;
  assign n11211 = n10772 ^ n3397;
  assign n11212 = ~n10956 & ~n11211;
  assign n11213 = n11212 ^ n10601;
  assign n11214 = n11213 ^ n11209;
  assign n11215 = n11210 & n11214;
  assign n11216 = n11215 ^ n3177;
  assign n11217 = n11216 ^ n2980;
  assign n11218 = n10776 & ~n10956;
  assign n11219 = n11218 ^ n10778;
  assign n11220 = n11219 ^ n11216;
  assign n11221 = n11217 & ~n11220;
  assign n11222 = n11221 ^ n2980;
  assign n11223 = n11222 ^ n2782;
  assign n11224 = n10782 & ~n10956;
  assign n11225 = n11224 ^ n10784;
  assign n11226 = n11225 ^ n11222;
  assign n11227 = n11223 & n11226;
  assign n11228 = n11227 ^ n2782;
  assign n11229 = n11228 ^ n2583;
  assign n11230 = n10788 & ~n10956;
  assign n11231 = n11230 ^ n10790;
  assign n11232 = n11231 ^ n11228;
  assign n11233 = n11229 & ~n11232;
  assign n11234 = n11233 ^ n2583;
  assign n11235 = n11234 ^ n2374;
  assign n11236 = n10794 & ~n10956;
  assign n11237 = n11236 ^ n10796;
  assign n11238 = n11237 ^ n11234;
  assign n11239 = n11235 & n11238;
  assign n11240 = n11239 ^ n2374;
  assign n11241 = n11240 ^ n2194;
  assign n11242 = n10800 & ~n10956;
  assign n11243 = n11242 ^ n10803;
  assign n11244 = n11243 ^ n11240;
  assign n11245 = ~n11241 & ~n11244;
  assign n11246 = n11245 ^ n2194;
  assign n11247 = n11246 ^ n2011;
  assign n11248 = ~n10807 & ~n10956;
  assign n11249 = n11248 ^ n10810;
  assign n11250 = n11249 ^ n11246;
  assign n11251 = ~n11247 & ~n11250;
  assign n11252 = n11251 ^ n2011;
  assign n11253 = n11252 ^ n1804;
  assign n11254 = ~n10814 & ~n10956;
  assign n11255 = n11254 ^ n10816;
  assign n11256 = n11255 ^ n11252;
  assign n11257 = n11253 & ~n11256;
  assign n11258 = n11257 ^ n1804;
  assign n11259 = n11258 ^ n1621;
  assign n11260 = n10820 & ~n10956;
  assign n11261 = n11260 ^ n10822;
  assign n11262 = n11261 ^ n11258;
  assign n11263 = n11259 & n11262;
  assign n11264 = n11263 ^ n1621;
  assign n11265 = n11264 ^ n1458;
  assign n11266 = n10826 & ~n10956;
  assign n11267 = n11266 ^ n10828;
  assign n11268 = n11267 ^ n11264;
  assign n11269 = n11265 & ~n11268;
  assign n11270 = n11269 ^ n1458;
  assign n11271 = n11270 ^ n1299;
  assign n11272 = n10832 & ~n10956;
  assign n11273 = n11272 ^ n10834;
  assign n11274 = n11273 ^ n11270;
  assign n11275 = n11271 & n11274;
  assign n11276 = n11275 ^ n1299;
  assign n11277 = n11276 ^ n10969;
  assign n11278 = n10970 & ~n11277;
  assign n11279 = n11278 ^ n1158;
  assign n11280 = n11279 ^ n10965;
  assign n11281 = ~n10966 & n11280;
  assign n11282 = n11281 ^ n1027;
  assign n11283 = n11282 ^ n905;
  assign n11284 = n10844 & ~n10956;
  assign n11285 = n11284 ^ n10847;
  assign n11286 = n11285 ^ n11282;
  assign n11287 = n11283 & ~n11286;
  assign n11288 = n11287 ^ n905;
  assign n11289 = n11288 ^ n803;
  assign n11290 = n10851 & ~n10956;
  assign n11291 = n11290 ^ n10854;
  assign n11292 = n11291 ^ n11288;
  assign n11293 = n11289 & n11292;
  assign n11294 = n11293 ^ n803;
  assign n11295 = n11294 ^ n707;
  assign n11296 = n10858 & ~n10956;
  assign n11297 = n11296 ^ n10860;
  assign n11298 = n11297 ^ n11294;
  assign n11299 = ~n11295 & ~n11298;
  assign n11300 = n11299 ^ n707;
  assign n11301 = n11300 ^ n608;
  assign n11302 = ~n10864 & ~n10956;
  assign n11303 = n11302 ^ n10866;
  assign n11304 = n11303 ^ n11300;
  assign n11305 = ~n11301 & ~n11304;
  assign n11306 = n11305 ^ n608;
  assign n11307 = n11306 ^ n514;
  assign n11308 = ~n10870 & ~n10956;
  assign n11309 = n11308 ^ n10872;
  assign n11310 = n11309 ^ n11306;
  assign n11311 = n11307 & ~n11310;
  assign n11312 = n11311 ^ n514;
  assign n11313 = n11312 ^ n436;
  assign n11314 = n10876 & ~n10956;
  assign n11315 = n11314 ^ n10878;
  assign n11316 = n11315 ^ n11312;
  assign n11317 = n11313 & n11316;
  assign n11318 = n11317 ^ n436;
  assign n11319 = ~n10962 & ~n11318;
  assign n11320 = ~n363 & ~n10961;
  assign n11321 = n10888 & ~n10956;
  assign n11322 = n11321 ^ n10890;
  assign n11323 = ~n11320 & ~n11322;
  assign n11324 = ~n11319 & n11323;
  assign n11325 = ~n10962 & n11322;
  assign n11326 = n11320 ^ n11318;
  assign n11327 = n11318 ^ n300;
  assign n11328 = n11318 & n11327;
  assign n11329 = n11328 ^ n11318;
  assign n11330 = ~n11326 & n11329;
  assign n11331 = n11330 ^ n11328;
  assign n11332 = n11331 ^ n11318;
  assign n11333 = n11332 ^ n300;
  assign n11334 = n11325 & n11333;
  assign n11335 = n11334 ^ n300;
  assign n11336 = ~n11324 & ~n11335;
  assign n11337 = n11336 ^ n243;
  assign n11338 = n10893 ^ n300;
  assign n11339 = ~n10956 & n11338;
  assign n11340 = n11339 ^ n10590;
  assign n11341 = n11340 ^ n11336;
  assign n11342 = ~n11337 & n11341;
  assign n11343 = n11342 ^ n243;
  assign n11344 = n11343 ^ n210;
  assign n11345 = n10896 ^ n243;
  assign n11346 = ~n10956 & n11345;
  assign n11347 = n11346 ^ n10587;
  assign n11348 = n11347 ^ n11343;
  assign n11349 = n11344 & ~n11348;
  assign n11350 = n11349 ^ n210;
  assign n11351 = n11350 ^ n147;
  assign n11352 = n10900 & ~n10956;
  assign n11353 = n11352 ^ n10902;
  assign n11354 = n11353 ^ n11350;
  assign n11355 = ~n11351 & ~n11354;
  assign n11356 = n11355 ^ n147;
  assign n11357 = ~n10959 & n11356;
  assign n11358 = n10916 & ~n10956;
  assign n11359 = n11358 ^ n10918;
  assign n11360 = ~n133 & ~n11359;
  assign n11361 = n132 & n10958;
  assign n11362 = ~n11360 & ~n11361;
  assign n11363 = ~n11357 & n11362;
  assign n11364 = n133 & n10909;
  assign n11365 = n10918 ^ n10916;
  assign n11366 = n11365 ^ n10955;
  assign n11367 = n10955 ^ n10915;
  assign n11368 = n10955 ^ n10918;
  assign n11369 = n10955 & ~n11368;
  assign n11370 = n11369 ^ n10955;
  assign n11371 = ~n11367 & n11370;
  assign n11372 = n11371 ^ n11369;
  assign n11373 = n11372 ^ n10955;
  assign n11374 = n11373 ^ n10918;
  assign n11375 = n11366 & ~n11374;
  assign n11376 = n11375 ^ n11365;
  assign n11377 = n11364 & n11376;
  assign n11382 = n10910 & n10955;
  assign n11378 = n1292 & ~n10918;
  assign n11379 = n10955 & n11378;
  assign n11380 = n10915 & n11379;
  assign n11381 = ~n10909 & ~n11380;
  assign n11383 = n11382 ^ n11381;
  assign n11384 = n11382 ^ n133;
  assign n11385 = n11382 ^ n10921;
  assign n11386 = ~n11382 & n11385;
  assign n11387 = n11386 ^ n11382;
  assign n11388 = ~n11384 & ~n11387;
  assign n11389 = n11388 ^ n11386;
  assign n11390 = n11389 ^ n11382;
  assign n11391 = n11390 ^ n10921;
  assign n11392 = n11383 & n11391;
  assign n11393 = n11392 ^ n11381;
  assign n11394 = ~n11377 & ~n11393;
  assign n11395 = ~n11363 & n11394;
  assign n11396 = n11356 ^ n132;
  assign n11397 = ~n11395 & n11396;
  assign n11398 = n11397 ^ n10958;
  assign n11399 = ~n133 & n11398;
  assign n11400 = n11283 & ~n11395;
  assign n11401 = n11400 ^ n11285;
  assign n11402 = n11401 ^ n803;
  assign n11403 = n11279 ^ n1027;
  assign n11404 = ~n11395 & n11403;
  assign n11405 = n11404 ^ n10965;
  assign n11406 = n11405 ^ n905;
  assign n11407 = n11253 & ~n11395;
  assign n11408 = n11407 ^ n11255;
  assign n11409 = ~n1621 & ~n11408;
  assign n11410 = n11259 & ~n11395;
  assign n11411 = n11410 ^ n11261;
  assign n11412 = ~n1458 & n11411;
  assign n11413 = ~n11409 & ~n11412;
  assign n11414 = ~n11247 & ~n11395;
  assign n11415 = n11414 ^ n11249;
  assign n11416 = n11415 ^ n1804;
  assign n11417 = ~n11241 & ~n11395;
  assign n11418 = n11417 ^ n11243;
  assign n11419 = n11418 ^ n2011;
  assign n11420 = n11235 & ~n11395;
  assign n11421 = n11420 ^ n11237;
  assign n11422 = n11421 ^ n2194;
  assign n11423 = n11229 & ~n11395;
  assign n11424 = n11423 ^ n11231;
  assign n11425 = n11424 ^ n2374;
  assign n11426 = n11197 & ~n11395;
  assign n11427 = n11426 ^ n11199;
  assign n11428 = n11427 ^ n3397;
  assign n11429 = n11182 ^ n4133;
  assign n11430 = n11184 ^ n11182;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = n11431 ^ n4133;
  assign n11433 = n11432 ^ n3882;
  assign n11434 = ~n11395 & n11433;
  assign n11435 = n11434 ^ n11187;
  assign n11436 = n11435 ^ n3634;
  assign n11437 = ~n11136 & ~n11138;
  assign n11438 = n10982 & ~n11437;
  assign n11439 = ~n11140 & ~n11438;
  assign n11440 = n11439 ^ n5108;
  assign n11441 = ~n11395 & ~n11440;
  assign n11442 = n11441 ^ n11142;
  assign n11443 = n11442 ^ n4851;
  assign n11444 = ~n10981 & ~n11437;
  assign n11445 = n11444 ^ n5363;
  assign n11446 = ~n11395 & n11445;
  assign n11447 = n11446 ^ n10976;
  assign n11448 = n11447 ^ n5108;
  assign n11449 = n11131 & ~n11395;
  assign n11450 = n11449 ^ n11133;
  assign n11451 = n11450 ^ n5625;
  assign n11452 = n11125 & ~n11395;
  assign n11453 = n11452 ^ n11127;
  assign n11454 = n11453 ^ n5905;
  assign n11455 = x24 & ~x25;
  assign n11456 = ~n10956 & n11455;
  assign n11457 = n11022 ^ n10585;
  assign n11458 = n11053 ^ n11022;
  assign n11459 = n11457 & n11458;
  assign n11460 = n11459 ^ n11022;
  assign n11461 = ~n11456 & ~n11460;
  assign n11462 = n11461 ^ n10229;
  assign n11463 = n10620 ^ n10585;
  assign n11464 = ~n10956 & n11463;
  assign n11465 = n11464 ^ n10585;
  assign n11466 = n11465 ^ x26;
  assign n11467 = n11466 ^ n11461;
  assign n11468 = n11462 & ~n11467;
  assign n11469 = n11468 ^ n10229;
  assign n11470 = n11469 ^ n9867;
  assign n11471 = ~n11395 & n11470;
  assign n11472 = n11471 ^ n11019;
  assign n11473 = n11472 ^ n9502;
  assign n11474 = ~n11395 & n11462;
  assign n11475 = n11474 ^ n11466;
  assign n11476 = n11475 ^ n9867;
  assign n11477 = ~x20 & ~x21;
  assign n11478 = n10956 & n11477;
  assign n11479 = ~x22 & n11478;
  assign n11480 = n11479 ^ n10956;
  assign n11481 = n11395 ^ x23;
  assign n11482 = ~n11480 & n11481;
  assign n11483 = ~n10956 & n11477;
  assign n11484 = n11483 ^ x23;
  assign n11485 = n11484 ^ n11483;
  assign n11486 = n11483 ^ n11395;
  assign n11487 = n11486 ^ n11483;
  assign n11488 = ~n11485 & ~n11487;
  assign n11489 = n11488 ^ n11483;
  assign n11490 = x22 & n11489;
  assign n11491 = n11490 ^ n11483;
  assign n11492 = ~n11482 & ~n11491;
  assign n11493 = n11492 ^ n10585;
  assign n11494 = n11021 ^ n10956;
  assign n11495 = ~n11395 & ~n11494;
  assign n11496 = n11495 ^ n10956;
  assign n11497 = n11496 ^ x24;
  assign n11498 = n11497 ^ n11492;
  assign n11499 = ~n11493 & n11498;
  assign n11500 = n11499 ^ n10585;
  assign n11501 = n11500 ^ n10229;
  assign n11503 = n11457 ^ x24;
  assign n11504 = n11503 ^ n11457;
  assign n11505 = n11457 ^ n11022;
  assign n11506 = n11504 & ~n11505;
  assign n11507 = n11506 ^ n11457;
  assign n11508 = ~n10956 & n11507;
  assign n11509 = n11508 ^ n11457;
  assign n11502 = ~x24 & ~n10956;
  assign n11510 = n11509 ^ n11502;
  assign n11511 = n11021 ^ n10585;
  assign n11512 = n11511 ^ n11509;
  assign n11513 = n11509 ^ n11395;
  assign n11514 = ~n11509 & n11513;
  assign n11515 = n11514 ^ n11509;
  assign n11516 = n11512 & ~n11515;
  assign n11517 = n11516 ^ n11514;
  assign n11518 = n11517 ^ n11509;
  assign n11519 = n11518 ^ n11395;
  assign n11520 = n11510 & n11519;
  assign n11521 = n11520 ^ n11502;
  assign n11522 = n11521 ^ x25;
  assign n11523 = n11522 ^ n11500;
  assign n11524 = ~n11501 & n11523;
  assign n11525 = n11524 ^ n10229;
  assign n11526 = n11525 ^ n11475;
  assign n11527 = n11476 & ~n11526;
  assign n11528 = n11527 ^ n9867;
  assign n11529 = n11528 ^ n11472;
  assign n11530 = n11473 & ~n11529;
  assign n11531 = n11530 ^ n9502;
  assign n11532 = n11531 ^ n9129;
  assign n11533 = n11079 ^ n9502;
  assign n11534 = ~n11395 & n11533;
  assign n11535 = n11534 ^ n10996;
  assign n11536 = n11535 ^ n11531;
  assign n11537 = n11532 & n11536;
  assign n11538 = n11537 ^ n9129;
  assign n11539 = n11538 ^ n8769;
  assign n11540 = n11083 & ~n11395;
  assign n11541 = n11540 ^ n11085;
  assign n11542 = n11541 ^ n11538;
  assign n11543 = n11539 & ~n11542;
  assign n11544 = n11543 ^ n8769;
  assign n11545 = n11544 ^ n8422;
  assign n11546 = n11089 & ~n11395;
  assign n11547 = n11546 ^ n11091;
  assign n11548 = n11547 ^ n11544;
  assign n11549 = n11545 & n11548;
  assign n11550 = n11549 ^ n8422;
  assign n11551 = n11550 ^ n8083;
  assign n11552 = n11095 & ~n11395;
  assign n11553 = n11552 ^ n11097;
  assign n11554 = n11553 ^ n11550;
  assign n11555 = n11551 & ~n11554;
  assign n11556 = n11555 ^ n8083;
  assign n11557 = n11556 ^ n7777;
  assign n11558 = n11100 ^ n8083;
  assign n11559 = ~n11395 & n11558;
  assign n11560 = n11559 ^ n10993;
  assign n11561 = n11560 ^ n11556;
  assign n11562 = n11557 & n11561;
  assign n11563 = n11562 ^ n7777;
  assign n11564 = n11563 ^ n7463;
  assign n11565 = n11103 ^ n7777;
  assign n11566 = ~n11395 & n11565;
  assign n11567 = n11566 ^ n10990;
  assign n11568 = n11567 ^ n11563;
  assign n11569 = n11564 & ~n11568;
  assign n11570 = n11569 ^ n7463;
  assign n11571 = n11570 ^ n7135;
  assign n11572 = n11106 ^ n7463;
  assign n11573 = ~n11395 & n11572;
  assign n11574 = n11573 ^ n10987;
  assign n11575 = n11574 ^ n11570;
  assign n11576 = n11571 & n11575;
  assign n11577 = n11576 ^ n7135;
  assign n11578 = n11577 ^ n6802;
  assign n11579 = n11109 ^ n7135;
  assign n11580 = ~n11395 & n11579;
  assign n11581 = n11580 ^ n10984;
  assign n11582 = n11581 ^ n11577;
  assign n11583 = n11578 & ~n11582;
  assign n11584 = n11583 ^ n6802;
  assign n11585 = n11584 ^ n6479;
  assign n11586 = n11113 & ~n11395;
  assign n11587 = n11586 ^ n11115;
  assign n11588 = n11587 ^ n11584;
  assign n11589 = n11585 & n11588;
  assign n11590 = n11589 ^ n6479;
  assign n11591 = n11590 ^ n6181;
  assign n11592 = n11119 & ~n11395;
  assign n11593 = n11592 ^ n11121;
  assign n11594 = n11593 ^ n11590;
  assign n11595 = n11591 & ~n11594;
  assign n11596 = n11595 ^ n6181;
  assign n11597 = n11596 ^ n11453;
  assign n11598 = ~n11454 & n11597;
  assign n11599 = n11598 ^ n5905;
  assign n11600 = n11599 ^ n11450;
  assign n11601 = n11451 & ~n11600;
  assign n11602 = n11601 ^ n5625;
  assign n11603 = n11602 ^ n5363;
  assign n11604 = n11136 ^ n5625;
  assign n11605 = ~n11395 & n11604;
  assign n11606 = n11605 ^ n10980;
  assign n11607 = n11606 ^ n11602;
  assign n11608 = n11603 & n11607;
  assign n11609 = n11608 ^ n5363;
  assign n11610 = n11609 ^ n11447;
  assign n11611 = n11448 & ~n11610;
  assign n11612 = n11611 ^ n5108;
  assign n11613 = n11612 ^ n11442;
  assign n11614 = n11443 & ~n11613;
  assign n11615 = n11614 ^ n4851;
  assign n11616 = n11615 ^ n4606;
  assign n11617 = n11144 & ~n11438;
  assign n11618 = ~n11149 & ~n11617;
  assign n11619 = n11618 ^ n4851;
  assign n11620 = ~n11395 & n11619;
  assign n11621 = n11620 ^ n10972;
  assign n11622 = n11621 ^ n11615;
  assign n11623 = n11616 & ~n11622;
  assign n11624 = n11623 ^ n4606;
  assign n11625 = n11624 ^ n4362;
  assign n11626 = n11155 ^ n4606;
  assign n11627 = ~n11395 & n11626;
  assign n11628 = n11627 ^ n11163;
  assign n11629 = n11628 ^ n11624;
  assign n11630 = n11625 & n11629;
  assign n11631 = n11630 ^ n4362;
  assign n11632 = n11631 ^ n4133;
  assign n11633 = n11163 ^ n11155;
  assign n11634 = n11626 & n11633;
  assign n11635 = n11634 ^ n4606;
  assign n11636 = n11635 ^ n4362;
  assign n11637 = ~n11395 & n11636;
  assign n11638 = n11637 ^ n11159;
  assign n11639 = n11638 ^ n11631;
  assign n11640 = n11632 & ~n11639;
  assign n11641 = n11640 ^ n4133;
  assign n11642 = n11641 ^ n3882;
  assign n11643 = ~n11395 & ~n11429;
  assign n11644 = n11643 ^ n11184;
  assign n11645 = n11644 ^ n11641;
  assign n11646 = n11642 & n11645;
  assign n11647 = n11646 ^ n3882;
  assign n11648 = n11647 ^ n11435;
  assign n11649 = ~n11436 & ~n11648;
  assign n11650 = n11649 ^ n3634;
  assign n11651 = n11650 ^ n11427;
  assign n11652 = ~n11428 & ~n11651;
  assign n11653 = n11652 ^ n3397;
  assign n11654 = n11653 ^ n3177;
  assign n11655 = ~n11203 & ~n11395;
  assign n11656 = n11655 ^ n11206;
  assign n11657 = n11656 ^ n11653;
  assign n11658 = n11654 & ~n11657;
  assign n11659 = n11658 ^ n3177;
  assign n11660 = n11659 ^ n2980;
  assign n11661 = n11210 & ~n11395;
  assign n11662 = n11661 ^ n11213;
  assign n11663 = n11662 ^ n11659;
  assign n11664 = n11660 & n11663;
  assign n11665 = n11664 ^ n2980;
  assign n11666 = n11665 ^ n2782;
  assign n11667 = n11217 & ~n11395;
  assign n11668 = n11667 ^ n11219;
  assign n11669 = n11668 ^ n11665;
  assign n11670 = n11666 & ~n11669;
  assign n11671 = n11670 ^ n2782;
  assign n11672 = n11671 ^ n2583;
  assign n11673 = n11223 & ~n11395;
  assign n11674 = n11673 ^ n11225;
  assign n11675 = n11674 ^ n11671;
  assign n11676 = n11672 & n11675;
  assign n11677 = n11676 ^ n2583;
  assign n11678 = n11677 ^ n11424;
  assign n11679 = n11425 & ~n11678;
  assign n11680 = n11679 ^ n2374;
  assign n11681 = n11680 ^ n11421;
  assign n11682 = n11422 & n11681;
  assign n11683 = n11682 ^ n2194;
  assign n11684 = n11683 ^ n11418;
  assign n11685 = n11419 & n11684;
  assign n11686 = n11685 ^ n2011;
  assign n11687 = n11686 ^ n11415;
  assign n11688 = ~n11416 & n11687;
  assign n11689 = n11688 ^ n1804;
  assign n11690 = n11413 & n11689;
  assign n11691 = n11411 ^ n1458;
  assign n11692 = n1621 & n11408;
  assign n11693 = n11692 ^ n11411;
  assign n11694 = ~n11691 & n11693;
  assign n11695 = n11694 ^ n1458;
  assign n11696 = ~n11690 & ~n11695;
  assign n11697 = n11696 ^ n1299;
  assign n11698 = n11265 & ~n11395;
  assign n11699 = n11698 ^ n11267;
  assign n11700 = n11699 ^ n11696;
  assign n11701 = ~n11697 & n11700;
  assign n11702 = n11701 ^ n1299;
  assign n11703 = n11702 ^ n1158;
  assign n11704 = n11271 & ~n11395;
  assign n11705 = n11704 ^ n11273;
  assign n11706 = n11705 ^ n11702;
  assign n11707 = n11703 & n11706;
  assign n11708 = n11707 ^ n1158;
  assign n11709 = n11708 ^ n1027;
  assign n11710 = n11276 ^ n1158;
  assign n11711 = ~n11395 & n11710;
  assign n11712 = n11711 ^ n10969;
  assign n11713 = n11712 ^ n11708;
  assign n11714 = n11709 & ~n11713;
  assign n11715 = n11714 ^ n1027;
  assign n11716 = n11715 ^ n11405;
  assign n11717 = ~n11406 & n11716;
  assign n11718 = n11717 ^ n905;
  assign n11719 = n11718 ^ n11401;
  assign n11720 = n11402 & ~n11719;
  assign n11721 = n11720 ^ n803;
  assign n11722 = n11721 ^ n707;
  assign n11723 = n11289 & ~n11395;
  assign n11724 = n11723 ^ n11291;
  assign n11725 = n11724 ^ n11721;
  assign n11726 = ~n11722 & n11725;
  assign n11727 = n11726 ^ n707;
  assign n11728 = n11727 ^ n608;
  assign n11729 = ~n11295 & ~n11395;
  assign n11730 = n11729 ^ n11297;
  assign n11731 = n11730 ^ n11727;
  assign n11732 = ~n11728 & n11731;
  assign n11733 = n11732 ^ n608;
  assign n11734 = n11733 ^ n514;
  assign n11735 = ~n11301 & ~n11395;
  assign n11736 = n11735 ^ n11303;
  assign n11737 = n11736 ^ n11733;
  assign n11738 = n11734 & n11737;
  assign n11739 = n11738 ^ n514;
  assign n11740 = n11739 ^ n436;
  assign n11741 = n11307 & ~n11395;
  assign n11742 = n11741 ^ n11309;
  assign n11743 = n11742 ^ n11739;
  assign n11744 = n11740 & ~n11743;
  assign n11745 = n11744 ^ n436;
  assign n11746 = n11745 ^ n363;
  assign n11747 = n11313 & ~n11395;
  assign n11748 = n11747 ^ n11315;
  assign n11749 = n11748 ^ n11745;
  assign n11750 = n11746 & n11749;
  assign n11751 = n11750 ^ n363;
  assign n11752 = n11751 ^ n300;
  assign n11753 = n11318 ^ n363;
  assign n11754 = ~n11395 & n11753;
  assign n11755 = n11754 ^ n10961;
  assign n11756 = n11755 ^ n11751;
  assign n11757 = n11752 & ~n11756;
  assign n11758 = n11757 ^ n300;
  assign n11759 = n11758 ^ n243;
  assign n11760 = ~n11319 & ~n11320;
  assign n11761 = n11760 ^ n300;
  assign n11762 = ~n11395 & n11761;
  assign n11763 = n11762 ^ n11322;
  assign n11764 = n11763 ^ n11758;
  assign n11765 = n11759 & n11764;
  assign n11766 = n11765 ^ n243;
  assign n11767 = n11766 ^ n210;
  assign n11768 = ~n11337 & ~n11395;
  assign n11769 = n11768 ^ n11340;
  assign n11770 = n11769 ^ n11766;
  assign n11771 = n11767 & ~n11770;
  assign n11772 = n11771 ^ n210;
  assign n11773 = n11772 ^ n147;
  assign n11774 = n11344 & ~n11395;
  assign n11775 = n11774 ^ n11347;
  assign n11776 = n11775 ^ n11772;
  assign n11777 = ~n11773 & ~n11776;
  assign n11778 = n11777 ^ n147;
  assign n11779 = n11778 ^ n132;
  assign n11780 = ~n11351 & ~n11395;
  assign n11781 = n11780 ^ n11353;
  assign n11782 = n11781 ^ n11778;
  assign n11783 = n11779 & n11782;
  assign n11784 = n11783 ^ n132;
  assign n11785 = ~n11399 & ~n11784;
  assign n11786 = ~n132 & ~n11356;
  assign n11787 = n11394 ^ n11359;
  assign n11788 = n133 & ~n11787;
  assign n11789 = n11788 ^ n11359;
  assign n11790 = ~n11786 & ~n11789;
  assign n11791 = n11359 ^ n11356;
  assign n11792 = ~n11396 & ~n11791;
  assign n11793 = n133 & n11792;
  assign n11794 = ~n11790 & ~n11793;
  assign n11795 = n10958 & ~n11794;
  assign n11796 = n1287 & ~n10958;
  assign n11797 = n11796 ^ n11356;
  assign n11798 = n11797 ^ n11796;
  assign n11799 = n1292 & ~n10958;
  assign n11800 = n11799 ^ n11796;
  assign n11801 = ~n11798 & n11800;
  assign n11802 = n11801 ^ n11796;
  assign n11803 = n132 & n11356;
  assign n11804 = n11803 ^ n11394;
  assign n11805 = n11394 ^ n133;
  assign n11806 = ~n11394 & n11805;
  assign n11807 = n11806 ^ n11394;
  assign n11808 = n11804 & ~n11807;
  assign n11809 = n11808 ^ n11806;
  assign n11810 = n11809 ^ n11394;
  assign n11811 = n11810 ^ n133;
  assign n11812 = ~n11802 & n11811;
  assign n11813 = n11812 ^ n11802;
  assign n11814 = ~n11359 & n11813;
  assign n11815 = ~n133 & n11359;
  assign n11816 = ~n11361 & n11815;
  assign n11817 = ~n11357 & n11816;
  assign n11818 = ~n11814 & ~n11817;
  assign n11819 = ~n11795 & n11818;
  assign n11820 = ~n11785 & ~n11819;
  assign n11821 = ~x16 & ~x17;
  assign n11822 = ~x18 & n11821;
  assign n11823 = n11820 & ~n11822;
  assign n11824 = n11767 & ~n11820;
  assign n11825 = n11824 ^ n11769;
  assign n11826 = n147 & ~n11825;
  assign n11827 = n11740 & ~n11820;
  assign n11828 = n11827 ^ n11742;
  assign n11829 = n11828 ^ n363;
  assign n11830 = n11734 & ~n11820;
  assign n11831 = n11830 ^ n11736;
  assign n11832 = n11831 ^ n436;
  assign n11833 = n11632 & ~n11820;
  assign n11834 = n11833 ^ n11638;
  assign n11835 = n11834 ^ n3882;
  assign n11836 = n11625 & ~n11820;
  assign n11837 = n11836 ^ n11628;
  assign n11838 = n11837 ^ n4133;
  assign n11839 = ~n11501 & ~n11820;
  assign n11840 = n11839 ^ n11522;
  assign n11841 = n11840 ^ n9867;
  assign n11842 = ~n11493 & ~n11820;
  assign n11843 = n11842 ^ n11497;
  assign n11844 = n11843 ^ n10229;
  assign n11846 = n11395 ^ n10956;
  assign n11847 = n11846 ^ n11395;
  assign n11848 = n11847 ^ n11846;
  assign n11849 = n11846 ^ n11477;
  assign n11850 = n11848 & n11849;
  assign n11851 = n11850 ^ n11846;
  assign n11852 = ~x22 & n11851;
  assign n11853 = n11852 ^ n11846;
  assign n11845 = ~x22 & ~n11395;
  assign n11854 = n11853 ^ n11845;
  assign n11855 = n11477 ^ n10956;
  assign n11856 = n11855 ^ n11853;
  assign n11857 = n11853 ^ n11820;
  assign n11858 = ~n11853 & n11857;
  assign n11859 = n11858 ^ n11853;
  assign n11860 = ~n11856 & ~n11859;
  assign n11861 = n11860 ^ n11858;
  assign n11862 = n11861 ^ n11853;
  assign n11863 = n11862 ^ n11820;
  assign n11864 = n11854 & n11863;
  assign n11865 = n11864 ^ n11845;
  assign n11866 = n11865 ^ x23;
  assign n11867 = n11866 ^ n10585;
  assign n11876 = x21 ^ x20;
  assign n11877 = n11876 ^ x20;
  assign n11869 = ~x18 & ~x19;
  assign n11870 = ~x20 & n11869;
  assign n11878 = n11395 & ~n11870;
  assign n11879 = n11878 ^ x20;
  assign n11880 = n11877 & ~n11879;
  assign n11881 = n11880 ^ x20;
  assign n11882 = n11881 ^ x21;
  assign n11883 = n11882 ^ n11881;
  assign n11884 = ~n11395 & n11870;
  assign n11885 = n11884 ^ n11881;
  assign n11886 = n11885 ^ n11881;
  assign n11887 = ~n11883 & n11886;
  assign n11888 = n11887 ^ n11881;
  assign n11889 = x22 & n11888;
  assign n11890 = n11889 ^ n11881;
  assign n11868 = n11395 ^ x22;
  assign n11871 = n11870 ^ n11395;
  assign n11872 = n11395 ^ x21;
  assign n11873 = ~n11871 & n11872;
  assign n11874 = n11873 ^ n11395;
  assign n11875 = n11868 & ~n11874;
  assign n11891 = n11890 ^ n11875;
  assign n11892 = n11820 & n11891;
  assign n11893 = n11892 ^ n11890;
  assign n11894 = ~x21 & n11820;
  assign n11895 = n11477 ^ n11395;
  assign n11896 = ~n11820 & ~n11895;
  assign n11897 = n11896 ^ n11395;
  assign n11898 = ~n11894 & ~n11897;
  assign n11899 = ~x22 & ~n11898;
  assign n11900 = x21 & ~n11820;
  assign n11901 = n11395 & ~n11900;
  assign n11902 = n11870 & ~n11901;
  assign n11903 = n11820 & ~n11870;
  assign n11904 = n11903 ^ x21;
  assign n11905 = n11903 ^ x22;
  assign n11906 = ~n11903 & ~n11905;
  assign n11907 = n11906 ^ n11903;
  assign n11908 = n11904 & ~n11907;
  assign n11909 = n11908 ^ n11906;
  assign n11910 = n11909 ^ n11903;
  assign n11911 = n11910 ^ x22;
  assign n11912 = n11395 & ~n11911;
  assign n11913 = n11912 ^ x22;
  assign n11914 = ~n11902 & ~n11913;
  assign n11915 = ~n11899 & n11914;
  assign n11916 = ~n10956 & ~n11915;
  assign n11917 = ~n11893 & ~n11916;
  assign n11918 = n11917 ^ n11866;
  assign n11919 = ~n11867 & ~n11918;
  assign n11920 = n11919 ^ n10585;
  assign n11921 = n11920 ^ n11843;
  assign n11922 = ~n11844 & ~n11921;
  assign n11923 = n11922 ^ n10229;
  assign n11924 = n11923 ^ n11840;
  assign n11925 = n11841 & ~n11924;
  assign n11926 = n11925 ^ n9867;
  assign n11927 = n11926 ^ n9502;
  assign n11928 = n11525 ^ n9867;
  assign n11929 = ~n11820 & n11928;
  assign n11930 = n11929 ^ n11475;
  assign n11931 = n11930 ^ n11926;
  assign n11932 = n11927 & ~n11931;
  assign n11933 = n11932 ^ n9502;
  assign n11934 = n11933 ^ n9129;
  assign n11935 = n11528 ^ n9502;
  assign n11936 = ~n11820 & n11935;
  assign n11937 = n11936 ^ n11472;
  assign n11938 = n11937 ^ n11933;
  assign n11939 = n11934 & ~n11938;
  assign n11940 = n11939 ^ n9129;
  assign n11941 = n11940 ^ n8769;
  assign n11942 = n11532 & ~n11820;
  assign n11943 = n11942 ^ n11535;
  assign n11944 = n11943 ^ n11940;
  assign n11945 = n11941 & n11944;
  assign n11946 = n11945 ^ n8769;
  assign n11947 = n11946 ^ n8422;
  assign n11948 = n11539 & ~n11820;
  assign n11949 = n11948 ^ n11541;
  assign n11950 = n11949 ^ n11946;
  assign n11951 = n11947 & ~n11950;
  assign n11952 = n11951 ^ n8422;
  assign n11953 = n11952 ^ n8083;
  assign n11954 = n11545 & ~n11820;
  assign n11955 = n11954 ^ n11547;
  assign n11956 = n11955 ^ n11952;
  assign n11957 = n11953 & n11956;
  assign n11958 = n11957 ^ n8083;
  assign n11959 = n11958 ^ n7777;
  assign n11960 = n11551 & ~n11820;
  assign n11961 = n11960 ^ n11553;
  assign n11962 = n11961 ^ n11958;
  assign n11963 = n11959 & ~n11962;
  assign n11964 = n11963 ^ n7777;
  assign n11965 = n11964 ^ n7463;
  assign n11966 = n11557 & ~n11820;
  assign n11967 = n11966 ^ n11560;
  assign n11968 = n11967 ^ n11964;
  assign n11969 = n11965 & n11968;
  assign n11970 = n11969 ^ n7463;
  assign n11971 = n11970 ^ n7135;
  assign n11972 = n11564 & ~n11820;
  assign n11973 = n11972 ^ n11567;
  assign n11974 = n11973 ^ n11970;
  assign n11975 = n11971 & ~n11974;
  assign n11976 = n11975 ^ n7135;
  assign n11977 = n11976 ^ n6802;
  assign n11978 = n11571 & ~n11820;
  assign n11979 = n11978 ^ n11574;
  assign n11980 = n11979 ^ n11976;
  assign n11981 = n11977 & n11980;
  assign n11982 = n11981 ^ n6802;
  assign n11983 = n11982 ^ n6479;
  assign n11984 = n11578 & ~n11820;
  assign n11985 = n11984 ^ n11581;
  assign n11986 = n11985 ^ n11982;
  assign n11987 = n11983 & ~n11986;
  assign n11988 = n11987 ^ n6479;
  assign n11989 = n11988 ^ n6181;
  assign n11990 = n11585 & ~n11820;
  assign n11991 = n11990 ^ n11587;
  assign n11992 = n11991 ^ n11988;
  assign n11993 = n11989 & n11992;
  assign n11994 = n11993 ^ n6181;
  assign n11995 = n11994 ^ n5905;
  assign n11996 = n11591 & ~n11820;
  assign n11997 = n11996 ^ n11593;
  assign n11998 = n11997 ^ n11994;
  assign n11999 = n11995 & ~n11998;
  assign n12000 = n11999 ^ n5905;
  assign n12001 = n12000 ^ n5625;
  assign n12002 = n11596 ^ n5905;
  assign n12003 = ~n11820 & n12002;
  assign n12004 = n12003 ^ n11453;
  assign n12005 = n12004 ^ n12000;
  assign n12006 = n12001 & n12005;
  assign n12007 = n12006 ^ n5625;
  assign n12008 = n12007 ^ n5363;
  assign n12009 = n11599 ^ n5625;
  assign n12010 = ~n11820 & n12009;
  assign n12011 = n12010 ^ n11450;
  assign n12012 = n12011 ^ n12007;
  assign n12013 = n12008 & ~n12012;
  assign n12014 = n12013 ^ n5363;
  assign n12015 = n12014 ^ n5108;
  assign n12016 = n11603 & ~n11820;
  assign n12017 = n12016 ^ n11606;
  assign n12018 = n12017 ^ n12014;
  assign n12019 = n12015 & n12018;
  assign n12020 = n12019 ^ n5108;
  assign n12021 = n12020 ^ n4851;
  assign n12022 = n11609 ^ n5108;
  assign n12023 = ~n11820 & n12022;
  assign n12024 = n12023 ^ n11447;
  assign n12025 = n12024 ^ n12020;
  assign n12026 = n12021 & ~n12025;
  assign n12027 = n12026 ^ n4851;
  assign n12028 = n12027 ^ n4606;
  assign n12029 = n11612 ^ n4851;
  assign n12030 = ~n11820 & n12029;
  assign n12031 = n12030 ^ n11442;
  assign n12032 = n12031 ^ n12027;
  assign n12033 = n12028 & ~n12032;
  assign n12034 = n12033 ^ n4606;
  assign n12035 = n12034 ^ n4362;
  assign n12036 = n11616 & ~n11820;
  assign n12037 = n12036 ^ n11621;
  assign n12038 = n12037 ^ n12034;
  assign n12039 = n12035 & ~n12038;
  assign n12040 = n12039 ^ n4362;
  assign n12041 = n12040 ^ n11837;
  assign n12042 = ~n11838 & n12041;
  assign n12043 = n12042 ^ n4133;
  assign n12044 = n12043 ^ n11834;
  assign n12045 = n11835 & ~n12044;
  assign n12046 = n12045 ^ n3882;
  assign n12047 = n12046 ^ n3634;
  assign n12048 = n11642 & ~n11820;
  assign n12049 = n12048 ^ n11644;
  assign n12050 = n12049 ^ n12046;
  assign n12051 = ~n12047 & n12050;
  assign n12052 = n12051 ^ n3634;
  assign n12053 = n12052 ^ n3397;
  assign n12054 = n11647 ^ n3634;
  assign n12055 = ~n11820 & ~n12054;
  assign n12056 = n12055 ^ n11435;
  assign n12057 = n12056 ^ n12052;
  assign n12058 = ~n12053 & n12057;
  assign n12059 = n12058 ^ n3397;
  assign n12060 = n12059 ^ n3177;
  assign n12061 = n11650 ^ n3397;
  assign n12062 = ~n11820 & ~n12061;
  assign n12063 = n12062 ^ n11427;
  assign n12064 = n12063 ^ n12059;
  assign n12065 = n12060 & n12064;
  assign n12066 = n12065 ^ n3177;
  assign n12067 = n12066 ^ n2980;
  assign n12068 = n11654 & ~n11820;
  assign n12069 = n12068 ^ n11656;
  assign n12070 = n12069 ^ n12066;
  assign n12071 = n12067 & ~n12070;
  assign n12072 = n12071 ^ n2980;
  assign n12073 = n12072 ^ n2782;
  assign n12074 = n11660 & ~n11820;
  assign n12075 = n12074 ^ n11662;
  assign n12076 = n12075 ^ n12072;
  assign n12077 = n12073 & n12076;
  assign n12078 = n12077 ^ n2782;
  assign n12079 = n12078 ^ n2583;
  assign n12080 = n11666 & ~n11820;
  assign n12081 = n12080 ^ n11668;
  assign n12082 = n12081 ^ n12078;
  assign n12083 = n12079 & ~n12082;
  assign n12084 = n12083 ^ n2583;
  assign n12085 = n12084 ^ n2374;
  assign n12086 = n11672 & ~n11820;
  assign n12087 = n12086 ^ n11674;
  assign n12088 = n12087 ^ n12084;
  assign n12089 = n12085 & n12088;
  assign n12090 = n12089 ^ n2374;
  assign n12091 = n12090 ^ n2194;
  assign n12092 = n11677 ^ n2374;
  assign n12093 = ~n11820 & n12092;
  assign n12094 = n12093 ^ n11424;
  assign n12095 = n12094 ^ n12090;
  assign n12096 = ~n12091 & ~n12095;
  assign n12097 = n12096 ^ n2194;
  assign n12098 = n12097 ^ n2011;
  assign n12099 = n11680 ^ n2194;
  assign n12100 = ~n11820 & ~n12099;
  assign n12101 = n12100 ^ n11421;
  assign n12102 = n12101 ^ n12097;
  assign n12103 = ~n12098 & ~n12102;
  assign n12104 = n12103 ^ n2011;
  assign n12105 = n12104 ^ n1804;
  assign n12106 = n11683 ^ n2011;
  assign n12107 = ~n11820 & ~n12106;
  assign n12108 = n12107 ^ n11418;
  assign n12109 = n12108 ^ n12104;
  assign n12110 = n12105 & ~n12109;
  assign n12111 = n12110 ^ n1804;
  assign n12112 = n12111 ^ n1621;
  assign n12113 = n11686 ^ n1804;
  assign n12114 = ~n11820 & n12113;
  assign n12115 = n12114 ^ n11415;
  assign n12116 = n12115 ^ n12111;
  assign n12117 = n12112 & n12116;
  assign n12118 = n12117 ^ n1621;
  assign n12119 = n12118 ^ n1458;
  assign n12120 = n11689 ^ n1621;
  assign n12121 = ~n11820 & n12120;
  assign n12122 = n12121 ^ n11408;
  assign n12123 = n12122 ^ n12118;
  assign n12124 = n12119 & ~n12123;
  assign n12125 = n12124 ^ n1458;
  assign n12126 = n12125 ^ n1299;
  assign n12127 = n11689 ^ n11408;
  assign n12128 = n12120 & ~n12127;
  assign n12129 = n12128 ^ n1621;
  assign n12130 = n12129 ^ n1458;
  assign n12131 = ~n11820 & n12130;
  assign n12132 = n12131 ^ n11411;
  assign n12133 = n12132 ^ n12125;
  assign n12134 = n12126 & n12133;
  assign n12135 = n12134 ^ n1299;
  assign n12136 = n12135 ^ n1158;
  assign n12137 = ~n11697 & ~n11820;
  assign n12138 = n12137 ^ n11699;
  assign n12139 = n12138 ^ n12135;
  assign n12140 = n12136 & ~n12139;
  assign n12141 = n12140 ^ n1158;
  assign n12142 = n12141 ^ n1027;
  assign n12143 = n11703 & ~n11820;
  assign n12144 = n12143 ^ n11705;
  assign n12145 = n12144 ^ n12141;
  assign n12146 = n12142 & n12145;
  assign n12147 = n12146 ^ n1027;
  assign n12148 = n12147 ^ n905;
  assign n12149 = n11709 & ~n11820;
  assign n12150 = n12149 ^ n11712;
  assign n12151 = n12150 ^ n12147;
  assign n12152 = n12148 & ~n12151;
  assign n12153 = n12152 ^ n905;
  assign n12154 = n12153 ^ n803;
  assign n12155 = n11715 ^ n905;
  assign n12156 = ~n11820 & n12155;
  assign n12157 = n12156 ^ n11405;
  assign n12158 = n12157 ^ n12153;
  assign n12159 = n12154 & n12158;
  assign n12160 = n12159 ^ n803;
  assign n12161 = n12160 ^ n707;
  assign n12162 = n11718 ^ n803;
  assign n12163 = ~n11820 & n12162;
  assign n12164 = n12163 ^ n11401;
  assign n12165 = n12164 ^ n12160;
  assign n12166 = ~n12161 & ~n12165;
  assign n12167 = n12166 ^ n707;
  assign n12168 = n12167 ^ n608;
  assign n12169 = ~n11722 & ~n11820;
  assign n12170 = n12169 ^ n11724;
  assign n12171 = n12170 ^ n12167;
  assign n12172 = ~n12168 & ~n12171;
  assign n12173 = n12172 ^ n608;
  assign n12174 = n12173 ^ n514;
  assign n12175 = ~n11728 & ~n11820;
  assign n12176 = n12175 ^ n11730;
  assign n12177 = n12176 ^ n12173;
  assign n12178 = n12174 & ~n12177;
  assign n12179 = n12178 ^ n514;
  assign n12180 = n12179 ^ n11831;
  assign n12181 = ~n11832 & n12180;
  assign n12182 = n12181 ^ n436;
  assign n12183 = n12182 ^ n11828;
  assign n12184 = n11829 & ~n12183;
  assign n12185 = n12184 ^ n363;
  assign n12186 = n12185 ^ n300;
  assign n12187 = n11746 & ~n11820;
  assign n12188 = n12187 ^ n11748;
  assign n12189 = n12188 ^ n12185;
  assign n12190 = n12186 & n12189;
  assign n12191 = n12190 ^ n300;
  assign n12192 = n12191 ^ n243;
  assign n12193 = n11752 & ~n11820;
  assign n12194 = n12193 ^ n11755;
  assign n12195 = n12194 ^ n12191;
  assign n12196 = n12192 & ~n12195;
  assign n12197 = n12196 ^ n243;
  assign n12198 = n12197 ^ n210;
  assign n12199 = n11759 & ~n11820;
  assign n12200 = n12199 ^ n11763;
  assign n12201 = n12200 ^ n12197;
  assign n12202 = n12198 & n12201;
  assign n12203 = n12202 ^ n210;
  assign n12204 = ~n11826 & n12203;
  assign n12205 = ~n147 & n11825;
  assign n12206 = ~n12204 & ~n12205;
  assign n12207 = ~n11773 & ~n11820;
  assign n12208 = n12207 ^ n11775;
  assign n12209 = ~n12206 & n12208;
  assign n12210 = ~n12205 & ~n12208;
  assign n12211 = ~n12204 & n12210;
  assign n12212 = ~n132 & ~n12211;
  assign n12213 = ~n12209 & ~n12212;
  assign n12214 = n11779 & ~n11820;
  assign n12215 = n12214 ^ n11781;
  assign n12216 = ~n133 & ~n12215;
  assign n12217 = ~n12213 & ~n12216;
  assign n12218 = n11398 & ~n11819;
  assign n12223 = n11398 ^ n132;
  assign n12224 = n12223 ^ n11783;
  assign n12225 = n12218 & n12224;
  assign n12226 = n12225 ^ n12224;
  assign n12219 = n11784 ^ n11398;
  assign n12220 = n12218 & ~n12219;
  assign n12221 = n12220 ^ n12219;
  assign n12222 = ~n12215 & n12221;
  assign n12227 = n12226 ^ n12222;
  assign n12228 = ~n133 & ~n12227;
  assign n12229 = n12228 ^ n12222;
  assign n12230 = ~n12217 & n12229;
  assign n12231 = n12230 ^ x19;
  assign n12232 = ~n11823 & n12231;
  assign n12234 = ~n11820 & n11821;
  assign n12233 = ~x19 & ~n12230;
  assign n12235 = n12234 ^ n12233;
  assign n12236 = ~x18 & n12235;
  assign n12237 = n12236 ^ n12233;
  assign n12238 = ~n12232 & ~n12237;
  assign n12239 = n12238 ^ n11395;
  assign n12240 = n11869 ^ n11820;
  assign n12241 = ~n12230 & ~n12240;
  assign n12242 = n12241 ^ n11820;
  assign n12243 = n12242 ^ x20;
  assign n12244 = n12243 ^ n12238;
  assign n12245 = n12239 & n12244;
  assign n12246 = n12245 ^ n11395;
  assign n12247 = n12246 ^ n10956;
  assign n12248 = n12192 & ~n12230;
  assign n12249 = n12248 ^ n12194;
  assign n12250 = n210 & n12249;
  assign n12251 = n12198 & ~n12230;
  assign n12252 = n12251 ^ n12200;
  assign n12253 = ~n147 & ~n12252;
  assign n12254 = ~n12250 & ~n12253;
  assign n12255 = n12182 ^ n363;
  assign n12256 = ~n12230 & n12255;
  assign n12257 = n12256 ^ n11828;
  assign n12258 = n12257 ^ n300;
  assign n12259 = n12179 ^ n436;
  assign n12260 = ~n12230 & n12259;
  assign n12261 = n12260 ^ n11831;
  assign n12262 = n12261 ^ n363;
  assign n12263 = n12174 & ~n12230;
  assign n12264 = n12263 ^ n12176;
  assign n12265 = n436 & n12264;
  assign n12266 = n12265 ^ n12261;
  assign n12267 = ~n12262 & ~n12266;
  assign n12268 = n12267 ^ n12261;
  assign n12269 = n12268 ^ n12257;
  assign n12270 = n12269 ^ n12257;
  assign n12271 = ~n12168 & ~n12230;
  assign n12272 = n12271 ^ n12170;
  assign n12273 = n514 & ~n12272;
  assign n12274 = n12085 & ~n12230;
  assign n12275 = n12274 ^ n12087;
  assign n12276 = n12275 ^ n2194;
  assign n12277 = n12079 & ~n12230;
  assign n12278 = n12277 ^ n12081;
  assign n12279 = n12278 ^ n2374;
  assign n12280 = n12043 ^ n3882;
  assign n12281 = ~n12230 & n12280;
  assign n12282 = n12281 ^ n11834;
  assign n12283 = n12282 ^ n3634;
  assign n12284 = n12040 ^ n4133;
  assign n12285 = ~n12230 & n12284;
  assign n12286 = n12285 ^ n11837;
  assign n12287 = n12286 ^ n3882;
  assign n12288 = n12021 & ~n12230;
  assign n12289 = n12288 ^ n12024;
  assign n12290 = n12289 ^ n4606;
  assign n12291 = n12015 & ~n12230;
  assign n12292 = n12291 ^ n12017;
  assign n12293 = n12292 ^ n4851;
  assign n12294 = n11995 & ~n12230;
  assign n12295 = n12294 ^ n11997;
  assign n12296 = n12295 ^ n5625;
  assign n12297 = n11989 & ~n12230;
  assign n12298 = n12297 ^ n11991;
  assign n12299 = n12298 ^ n5905;
  assign n12300 = n11920 ^ n10229;
  assign n12301 = ~n12230 & ~n12300;
  assign n12302 = n12301 ^ n11843;
  assign n12303 = n12302 ^ n9867;
  assign n12304 = n11917 ^ n10585;
  assign n12305 = ~n12230 & ~n12304;
  assign n12306 = n12305 ^ n11866;
  assign n12307 = n12306 ^ n10229;
  assign n12308 = n11903 ^ n11395;
  assign n12309 = ~x20 & ~n11820;
  assign n12310 = ~n11903 & n12309;
  assign n12311 = n12308 & n12310;
  assign n12312 = n12311 ^ n12308;
  assign n12313 = n12312 ^ n12309;
  assign n12314 = n11869 ^ n11395;
  assign n12315 = n12314 ^ n12312;
  assign n12316 = n12312 ^ n12230;
  assign n12317 = ~n12312 & n12316;
  assign n12318 = n12317 ^ n12312;
  assign n12319 = ~n12315 & ~n12318;
  assign n12320 = n12319 ^ n12317;
  assign n12321 = n12320 ^ n12312;
  assign n12322 = n12321 ^ n12230;
  assign n12323 = n12313 & n12322;
  assign n12324 = n12323 ^ n12309;
  assign n12325 = n12324 ^ x21;
  assign n12326 = n12325 ^ n12246;
  assign n12327 = n12247 & ~n12326;
  assign n12328 = n12327 ^ n10956;
  assign n12329 = n12328 ^ n10585;
  assign n12339 = n11897 ^ x22;
  assign n12330 = x20 & ~x21;
  assign n12331 = ~n11820 & n12330;
  assign n12332 = n11820 ^ x21;
  assign n12333 = n12332 ^ n11870;
  assign n12334 = ~n11871 & n12333;
  assign n12335 = n12334 ^ n11870;
  assign n12336 = ~n12331 & ~n12335;
  assign n12337 = n12336 ^ n10956;
  assign n12338 = ~n12230 & n12337;
  assign n12340 = n12339 ^ n12338;
  assign n12341 = n12340 ^ n12328;
  assign n12342 = ~n12329 & n12341;
  assign n12343 = n12342 ^ n10585;
  assign n12344 = n12343 ^ n12306;
  assign n12345 = n12307 & n12344;
  assign n12346 = n12345 ^ n10229;
  assign n12347 = n12346 ^ n12302;
  assign n12348 = ~n12303 & n12347;
  assign n12349 = n12348 ^ n9867;
  assign n12350 = n12349 ^ n9502;
  assign n12351 = n11923 ^ n9867;
  assign n12352 = ~n12230 & n12351;
  assign n12353 = n12352 ^ n11840;
  assign n12354 = n12353 ^ n12349;
  assign n12355 = n12350 & ~n12354;
  assign n12356 = n12355 ^ n9502;
  assign n12357 = n12356 ^ n9129;
  assign n12358 = n11927 & ~n12230;
  assign n12359 = n12358 ^ n11930;
  assign n12360 = n12359 ^ n12356;
  assign n12361 = n12357 & ~n12360;
  assign n12362 = n12361 ^ n9129;
  assign n12363 = n12362 ^ n8769;
  assign n12364 = n11934 & ~n12230;
  assign n12365 = n12364 ^ n11937;
  assign n12366 = n12365 ^ n12362;
  assign n12367 = n12363 & ~n12366;
  assign n12368 = n12367 ^ n8769;
  assign n12369 = n12368 ^ n8422;
  assign n12370 = n11941 & ~n12230;
  assign n12371 = n12370 ^ n11943;
  assign n12372 = n12371 ^ n12368;
  assign n12373 = n12369 & n12372;
  assign n12374 = n12373 ^ n8422;
  assign n12375 = n12374 ^ n8083;
  assign n12376 = n11947 & ~n12230;
  assign n12377 = n12376 ^ n11949;
  assign n12378 = n12377 ^ n12374;
  assign n12379 = n12375 & ~n12378;
  assign n12380 = n12379 ^ n8083;
  assign n12381 = n12380 ^ n7777;
  assign n12382 = n11953 & ~n12230;
  assign n12383 = n12382 ^ n11955;
  assign n12384 = n12383 ^ n12380;
  assign n12385 = n12381 & n12384;
  assign n12386 = n12385 ^ n7777;
  assign n12387 = n12386 ^ n7463;
  assign n12388 = n11959 & ~n12230;
  assign n12389 = n12388 ^ n11961;
  assign n12390 = n12389 ^ n12386;
  assign n12391 = n12387 & ~n12390;
  assign n12392 = n12391 ^ n7463;
  assign n12393 = n12392 ^ n7135;
  assign n12394 = n11965 & ~n12230;
  assign n12395 = n12394 ^ n11967;
  assign n12396 = n12395 ^ n12392;
  assign n12397 = n12393 & n12396;
  assign n12398 = n12397 ^ n7135;
  assign n12399 = n12398 ^ n6802;
  assign n12400 = n11971 & ~n12230;
  assign n12401 = n12400 ^ n11973;
  assign n12402 = n12401 ^ n12398;
  assign n12403 = n12399 & ~n12402;
  assign n12404 = n12403 ^ n6802;
  assign n12405 = n12404 ^ n6479;
  assign n12406 = n11977 & ~n12230;
  assign n12407 = n12406 ^ n11979;
  assign n12408 = n12407 ^ n12404;
  assign n12409 = n12405 & n12408;
  assign n12410 = n12409 ^ n6479;
  assign n12411 = n12410 ^ n6181;
  assign n12412 = n11983 & ~n12230;
  assign n12413 = n12412 ^ n11985;
  assign n12414 = n12413 ^ n12410;
  assign n12415 = n12411 & ~n12414;
  assign n12416 = n12415 ^ n6181;
  assign n12417 = n12416 ^ n12298;
  assign n12418 = ~n12299 & n12417;
  assign n12419 = n12418 ^ n5905;
  assign n12420 = n12419 ^ n12295;
  assign n12421 = n12296 & ~n12420;
  assign n12422 = n12421 ^ n5625;
  assign n12423 = n12422 ^ n5363;
  assign n12424 = n12001 & ~n12230;
  assign n12425 = n12424 ^ n12004;
  assign n12426 = n12425 ^ n12422;
  assign n12427 = n12423 & n12426;
  assign n12428 = n12427 ^ n5363;
  assign n12429 = n12428 ^ n5108;
  assign n12430 = n12008 & ~n12230;
  assign n12431 = n12430 ^ n12011;
  assign n12432 = n12431 ^ n12428;
  assign n12433 = n12429 & ~n12432;
  assign n12434 = n12433 ^ n5108;
  assign n12435 = n12434 ^ n12292;
  assign n12436 = ~n12293 & n12435;
  assign n12437 = n12436 ^ n4851;
  assign n12438 = n12437 ^ n12289;
  assign n12439 = n12290 & ~n12438;
  assign n12440 = n12439 ^ n4606;
  assign n12441 = n12440 ^ n4362;
  assign n12442 = n12028 & ~n12230;
  assign n12443 = n12442 ^ n12031;
  assign n12444 = n12443 ^ n12440;
  assign n12445 = n12441 & ~n12444;
  assign n12446 = n12445 ^ n4362;
  assign n12447 = n12446 ^ n4133;
  assign n12448 = n12035 & ~n12230;
  assign n12449 = n12448 ^ n12037;
  assign n12450 = n12449 ^ n12446;
  assign n12451 = n12447 & ~n12450;
  assign n12452 = n12451 ^ n4133;
  assign n12453 = n12452 ^ n12286;
  assign n12454 = ~n12287 & n12453;
  assign n12455 = n12454 ^ n3882;
  assign n12456 = n12455 ^ n12282;
  assign n12457 = ~n12283 & ~n12456;
  assign n12458 = n12457 ^ n3634;
  assign n12459 = n12458 ^ n3397;
  assign n12460 = ~n12047 & ~n12230;
  assign n12461 = n12460 ^ n12049;
  assign n12462 = n12461 ^ n12458;
  assign n12463 = ~n12459 & ~n12462;
  assign n12464 = n12463 ^ n3397;
  assign n12465 = n12464 ^ n3177;
  assign n12466 = ~n12053 & ~n12230;
  assign n12467 = n12466 ^ n12056;
  assign n12468 = n12467 ^ n12464;
  assign n12469 = n12465 & ~n12468;
  assign n12470 = n12469 ^ n3177;
  assign n12471 = n12470 ^ n2980;
  assign n12472 = n12060 & ~n12230;
  assign n12473 = n12472 ^ n12063;
  assign n12474 = n12473 ^ n12470;
  assign n12475 = n12471 & n12474;
  assign n12476 = n12475 ^ n2980;
  assign n12477 = n12476 ^ n2782;
  assign n12478 = n12067 & ~n12230;
  assign n12479 = n12478 ^ n12069;
  assign n12480 = n12479 ^ n12476;
  assign n12481 = n12477 & ~n12480;
  assign n12482 = n12481 ^ n2782;
  assign n12483 = n12482 ^ n2583;
  assign n12484 = n12073 & ~n12230;
  assign n12485 = n12484 ^ n12075;
  assign n12486 = n12485 ^ n12482;
  assign n12487 = n12483 & n12486;
  assign n12488 = n12487 ^ n2583;
  assign n12489 = n12488 ^ n12278;
  assign n12490 = n12279 & ~n12489;
  assign n12491 = n12490 ^ n2374;
  assign n12492 = n12491 ^ n12275;
  assign n12493 = n12276 & n12492;
  assign n12494 = n12493 ^ n2194;
  assign n12495 = n12494 ^ n2011;
  assign n12496 = ~n12091 & ~n12230;
  assign n12497 = n12496 ^ n12094;
  assign n12498 = n12497 ^ n12494;
  assign n12499 = ~n12495 & n12498;
  assign n12500 = n12499 ^ n2011;
  assign n12501 = n12500 ^ n1804;
  assign n12502 = ~n12098 & ~n12230;
  assign n12503 = n12502 ^ n12101;
  assign n12504 = n12503 ^ n12500;
  assign n12505 = n12501 & n12504;
  assign n12506 = n12505 ^ n1804;
  assign n12507 = n12506 ^ n1621;
  assign n12508 = n12105 & ~n12230;
  assign n12509 = n12508 ^ n12108;
  assign n12510 = n12509 ^ n12506;
  assign n12511 = n12507 & ~n12510;
  assign n12512 = n12511 ^ n1621;
  assign n12513 = n12512 ^ n1458;
  assign n12514 = n12112 & ~n12230;
  assign n12515 = n12514 ^ n12115;
  assign n12516 = n12515 ^ n12512;
  assign n12517 = n12513 & n12516;
  assign n12518 = n12517 ^ n1458;
  assign n12519 = n12518 ^ n1299;
  assign n12520 = n12119 & ~n12230;
  assign n12521 = n12520 ^ n12122;
  assign n12522 = n12521 ^ n12518;
  assign n12523 = n12519 & ~n12522;
  assign n12524 = n12523 ^ n1299;
  assign n12525 = n12524 ^ n1158;
  assign n12526 = n12126 & ~n12230;
  assign n12527 = n12526 ^ n12132;
  assign n12528 = n12527 ^ n12524;
  assign n12529 = n12525 & n12528;
  assign n12530 = n12529 ^ n1158;
  assign n12531 = n12530 ^ n1027;
  assign n12532 = n12136 & ~n12230;
  assign n12533 = n12532 ^ n12138;
  assign n12534 = n12533 ^ n12530;
  assign n12535 = n12531 & ~n12534;
  assign n12536 = n12535 ^ n1027;
  assign n12537 = n12536 ^ n905;
  assign n12538 = n12142 & ~n12230;
  assign n12539 = n12538 ^ n12144;
  assign n12540 = n12539 ^ n12536;
  assign n12541 = n12537 & n12540;
  assign n12542 = n12541 ^ n905;
  assign n12543 = n12542 ^ n803;
  assign n12544 = n12148 & ~n12230;
  assign n12545 = n12544 ^ n12150;
  assign n12546 = n12545 ^ n12542;
  assign n12547 = n12543 & ~n12546;
  assign n12548 = n12547 ^ n803;
  assign n12549 = n12548 ^ n707;
  assign n12550 = n12154 & ~n12230;
  assign n12551 = n12550 ^ n12157;
  assign n12552 = n12551 ^ n12548;
  assign n12553 = ~n12549 & n12552;
  assign n12554 = n12553 ^ n707;
  assign n12555 = n12554 ^ n608;
  assign n12556 = ~n12161 & ~n12230;
  assign n12557 = n12556 ^ n12164;
  assign n12558 = n12557 ^ n12554;
  assign n12559 = ~n12555 & n12558;
  assign n12560 = n12559 ^ n608;
  assign n12561 = ~n12273 & ~n12560;
  assign n12562 = ~n436 & ~n12264;
  assign n12563 = ~n514 & n12272;
  assign n12564 = ~n12562 & ~n12563;
  assign n12565 = ~n363 & n12261;
  assign n12566 = n12564 & ~n12565;
  assign n12567 = ~n12561 & n12566;
  assign n12568 = n12567 ^ n12257;
  assign n12569 = n12568 ^ n12257;
  assign n12570 = n12270 & ~n12569;
  assign n12571 = n12570 ^ n12257;
  assign n12572 = n12258 & n12571;
  assign n12573 = n12572 ^ n300;
  assign n12574 = n12573 ^ n243;
  assign n12575 = n12186 & ~n12230;
  assign n12576 = n12575 ^ n12188;
  assign n12577 = n12576 ^ n12573;
  assign n12578 = n12574 & n12577;
  assign n12579 = n12578 ^ n243;
  assign n12580 = n12254 & ~n12579;
  assign n12581 = n12203 ^ n147;
  assign n12582 = ~n12230 & ~n12581;
  assign n12583 = n12582 ^ n11825;
  assign n12584 = n12252 ^ n147;
  assign n12585 = ~n210 & ~n12249;
  assign n12586 = n12585 ^ n12252;
  assign n12587 = n12584 & ~n12586;
  assign n12588 = n12587 ^ n147;
  assign n12589 = n12583 & ~n12588;
  assign n12590 = ~n12580 & n12589;
  assign n12591 = n132 & ~n12590;
  assign n12592 = ~n12580 & ~n12588;
  assign n12593 = ~n12583 & ~n12592;
  assign n12594 = ~n12591 & ~n12593;
  assign n12595 = n12206 ^ n132;
  assign n12596 = ~n12230 & n12595;
  assign n12597 = n12596 ^ n12208;
  assign n12598 = ~n133 & ~n12597;
  assign n12599 = n12594 & ~n12598;
  assign n12600 = ~n12208 & n12229;
  assign n12601 = ~n12215 & ~n12600;
  assign n12602 = n12226 ^ n133;
  assign n12603 = n12602 ^ n12226;
  assign n12604 = ~n132 & n12209;
  assign n12605 = n12604 ^ n12226;
  assign n12606 = n12603 & ~n12605;
  assign n12607 = n12606 ^ n12226;
  assign n12608 = ~n12213 & n12607;
  assign n12609 = n12608 ^ n133;
  assign n12610 = n12601 & n12609;
  assign n12611 = ~n133 & ~n12213;
  assign n12612 = n12211 & n12215;
  assign n12613 = n1292 & n12612;
  assign n12614 = n12613 ^ n12215;
  assign n12615 = ~n12611 & n12614;
  assign n12616 = ~n12610 & ~n12615;
  assign n12617 = ~n12599 & n12616;
  assign n12618 = n12247 & ~n12617;
  assign n12619 = n12618 ^ n12325;
  assign n12620 = n12619 ^ n10585;
  assign n12621 = n12239 & ~n12617;
  assign n12622 = n12621 ^ n12243;
  assign n12623 = n12622 ^ n10956;
  assign n12624 = ~x14 & ~x15;
  assign n12625 = ~x16 & n12624;
  assign n12626 = n12230 & ~n12625;
  assign n12627 = n12617 ^ x17;
  assign n12628 = ~n12626 & n12627;
  assign n12630 = ~n12230 & n12624;
  assign n12629 = ~x17 & ~n12617;
  assign n12631 = n12630 ^ n12629;
  assign n12632 = ~x16 & n12631;
  assign n12633 = n12632 ^ n12629;
  assign n12634 = ~n12628 & ~n12633;
  assign n12635 = n12634 ^ n11820;
  assign n12638 = n11821 ^ x18;
  assign n12636 = n12230 ^ n11821;
  assign n12637 = n12617 & ~n12636;
  assign n12639 = n12638 ^ n12637;
  assign n12640 = n12639 ^ n12634;
  assign n12641 = n12635 & ~n12640;
  assign n12642 = n12641 ^ n11820;
  assign n12643 = n12642 ^ n11395;
  assign n12645 = n11822 ^ n11820;
  assign n12646 = n12645 ^ x18;
  assign n12647 = n12646 ^ n12645;
  assign n12648 = n12645 ^ n11822;
  assign n12649 = n12647 & n12648;
  assign n12650 = n12649 ^ n12645;
  assign n12651 = ~n12230 & ~n12650;
  assign n12652 = n12651 ^ n12645;
  assign n12644 = ~x18 & ~n12230;
  assign n12653 = n12652 ^ n12644;
  assign n12654 = n11821 ^ n11820;
  assign n12655 = n12654 ^ n12652;
  assign n12656 = n12652 ^ n12617;
  assign n12657 = n12652 & ~n12656;
  assign n12658 = n12657 ^ n12652;
  assign n12659 = n12655 & n12658;
  assign n12660 = n12659 ^ n12657;
  assign n12661 = n12660 ^ n12652;
  assign n12662 = n12661 ^ n12617;
  assign n12663 = ~n12653 & ~n12662;
  assign n12664 = n12663 ^ n12644;
  assign n12665 = n12664 ^ x19;
  assign n12666 = n12665 ^ n12642;
  assign n12667 = n12643 & ~n12666;
  assign n12668 = n12667 ^ n11395;
  assign n12669 = n12668 ^ n12622;
  assign n12670 = ~n12623 & n12669;
  assign n12671 = n12670 ^ n10956;
  assign n12672 = n12671 ^ n12619;
  assign n12673 = ~n12620 & ~n12672;
  assign n12674 = n12673 ^ n10585;
  assign n12675 = n12674 ^ n10229;
  assign n12676 = ~n12329 & ~n12617;
  assign n12677 = n12676 ^ n12340;
  assign n12678 = n12677 ^ n12674;
  assign n12679 = ~n12675 & ~n12678;
  assign n12680 = n12679 ^ n10229;
  assign n12681 = n12680 ^ n9867;
  assign n12682 = n12579 ^ n210;
  assign n12683 = ~n12617 & n12682;
  assign n12684 = n12683 ^ n12249;
  assign n12685 = n12684 ^ n147;
  assign n12686 = n12574 & ~n12617;
  assign n12687 = n12686 ^ n12576;
  assign n12688 = n12687 ^ n210;
  assign n12689 = n12491 ^ n2194;
  assign n12690 = ~n12617 & ~n12689;
  assign n12691 = n12690 ^ n12275;
  assign n12692 = n12691 ^ n2011;
  assign n12693 = n12488 ^ n2374;
  assign n12694 = ~n12617 & n12693;
  assign n12695 = n12694 ^ n12278;
  assign n12696 = n12695 ^ n2194;
  assign n12697 = n12369 & ~n12617;
  assign n12698 = n12697 ^ n12371;
  assign n12699 = n12698 ^ n8083;
  assign n12700 = n12363 & ~n12617;
  assign n12701 = n12700 ^ n12365;
  assign n12702 = n12701 ^ n8422;
  assign n12703 = n12343 ^ n10229;
  assign n12704 = ~n12617 & ~n12703;
  assign n12705 = n12704 ^ n12306;
  assign n12706 = n12705 ^ n12680;
  assign n12707 = n12681 & ~n12706;
  assign n12708 = n12707 ^ n9867;
  assign n12709 = n12708 ^ n9502;
  assign n12710 = n12346 ^ n9867;
  assign n12711 = ~n12617 & n12710;
  assign n12712 = n12711 ^ n12302;
  assign n12713 = n12712 ^ n12708;
  assign n12714 = n12709 & n12713;
  assign n12715 = n12714 ^ n9502;
  assign n12716 = n12715 ^ n9129;
  assign n12717 = n12350 & ~n12617;
  assign n12718 = n12717 ^ n12353;
  assign n12719 = n12718 ^ n12715;
  assign n12720 = n12716 & ~n12719;
  assign n12721 = n12720 ^ n9129;
  assign n12722 = n12721 ^ n8769;
  assign n12723 = n12357 & ~n12617;
  assign n12724 = n12723 ^ n12359;
  assign n12725 = n12724 ^ n12721;
  assign n12726 = n12722 & ~n12725;
  assign n12727 = n12726 ^ n8769;
  assign n12728 = n12727 ^ n12701;
  assign n12729 = n12702 & ~n12728;
  assign n12730 = n12729 ^ n8422;
  assign n12731 = n12730 ^ n12698;
  assign n12732 = ~n12699 & n12731;
  assign n12733 = n12732 ^ n8083;
  assign n12734 = n12733 ^ n7777;
  assign n12735 = n12375 & ~n12617;
  assign n12736 = n12735 ^ n12377;
  assign n12737 = n12736 ^ n12733;
  assign n12738 = n12734 & ~n12737;
  assign n12739 = n12738 ^ n7777;
  assign n12740 = n12739 ^ n7463;
  assign n12741 = n12381 & ~n12617;
  assign n12742 = n12741 ^ n12383;
  assign n12743 = n12742 ^ n12739;
  assign n12744 = n12740 & n12743;
  assign n12745 = n12744 ^ n7463;
  assign n12746 = n12745 ^ n7135;
  assign n12747 = n12387 & ~n12617;
  assign n12748 = n12747 ^ n12389;
  assign n12749 = n12748 ^ n12745;
  assign n12750 = n12746 & ~n12749;
  assign n12751 = n12750 ^ n7135;
  assign n12752 = n12751 ^ n6802;
  assign n12753 = n12393 & ~n12617;
  assign n12754 = n12753 ^ n12395;
  assign n12755 = n12754 ^ n12751;
  assign n12756 = n12752 & n12755;
  assign n12757 = n12756 ^ n6802;
  assign n12758 = n12757 ^ n6479;
  assign n12759 = n12399 & ~n12617;
  assign n12760 = n12759 ^ n12401;
  assign n12761 = n12760 ^ n12757;
  assign n12762 = n12758 & ~n12761;
  assign n12763 = n12762 ^ n6479;
  assign n12764 = n12763 ^ n6181;
  assign n12765 = n12405 & ~n12617;
  assign n12766 = n12765 ^ n12407;
  assign n12767 = n12766 ^ n12763;
  assign n12768 = n12764 & n12767;
  assign n12769 = n12768 ^ n6181;
  assign n12770 = n12769 ^ n5905;
  assign n12771 = n12411 & ~n12617;
  assign n12772 = n12771 ^ n12413;
  assign n12773 = n12772 ^ n12769;
  assign n12774 = n12770 & ~n12773;
  assign n12775 = n12774 ^ n5905;
  assign n12776 = n12775 ^ n5625;
  assign n12777 = n12416 ^ n5905;
  assign n12778 = ~n12617 & n12777;
  assign n12779 = n12778 ^ n12298;
  assign n12780 = n12779 ^ n12775;
  assign n12781 = n12776 & n12780;
  assign n12782 = n12781 ^ n5625;
  assign n12783 = n12782 ^ n5363;
  assign n12784 = n12419 ^ n5625;
  assign n12785 = ~n12617 & n12784;
  assign n12786 = n12785 ^ n12295;
  assign n12787 = n12786 ^ n12782;
  assign n12788 = n12783 & ~n12787;
  assign n12789 = n12788 ^ n5363;
  assign n12790 = n12789 ^ n5108;
  assign n12791 = n12423 & ~n12617;
  assign n12792 = n12791 ^ n12425;
  assign n12793 = n12792 ^ n12789;
  assign n12794 = n12790 & n12793;
  assign n12795 = n12794 ^ n5108;
  assign n12796 = n12795 ^ n4851;
  assign n12797 = n12429 & ~n12617;
  assign n12798 = n12797 ^ n12431;
  assign n12799 = n12798 ^ n12795;
  assign n12800 = n12796 & ~n12799;
  assign n12801 = n12800 ^ n4851;
  assign n12802 = n12801 ^ n4606;
  assign n12803 = n12434 ^ n4851;
  assign n12804 = ~n12617 & n12803;
  assign n12805 = n12804 ^ n12292;
  assign n12806 = n12805 ^ n12801;
  assign n12807 = n12802 & n12806;
  assign n12808 = n12807 ^ n4606;
  assign n12809 = n12808 ^ n4362;
  assign n12810 = n12437 ^ n4606;
  assign n12811 = ~n12617 & n12810;
  assign n12812 = n12811 ^ n12289;
  assign n12813 = n12812 ^ n12808;
  assign n12814 = n12809 & ~n12813;
  assign n12815 = n12814 ^ n4362;
  assign n12816 = n12815 ^ n4133;
  assign n12817 = n12441 & ~n12617;
  assign n12818 = n12817 ^ n12443;
  assign n12819 = n12818 ^ n12815;
  assign n12820 = n12816 & ~n12819;
  assign n12821 = n12820 ^ n4133;
  assign n12822 = n12821 ^ n3882;
  assign n12823 = n12447 & ~n12617;
  assign n12824 = n12823 ^ n12449;
  assign n12825 = n12824 ^ n12821;
  assign n12826 = n12822 & ~n12825;
  assign n12827 = n12826 ^ n3882;
  assign n12828 = n12827 ^ n3634;
  assign n12829 = n12452 ^ n3882;
  assign n12830 = ~n12617 & n12829;
  assign n12831 = n12830 ^ n12286;
  assign n12832 = n12831 ^ n12827;
  assign n12833 = ~n12828 & n12832;
  assign n12834 = n12833 ^ n3634;
  assign n12835 = n12834 ^ n3397;
  assign n12836 = n12455 ^ n3634;
  assign n12837 = ~n12617 & ~n12836;
  assign n12838 = n12837 ^ n12282;
  assign n12839 = n12838 ^ n12834;
  assign n12840 = ~n12835 & n12839;
  assign n12841 = n12840 ^ n3397;
  assign n12842 = n12841 ^ n3177;
  assign n12843 = ~n12459 & ~n12617;
  assign n12844 = n12843 ^ n12461;
  assign n12845 = n12844 ^ n12841;
  assign n12846 = n12842 & n12845;
  assign n12847 = n12846 ^ n3177;
  assign n12848 = n12847 ^ n2980;
  assign n12849 = n12465 & ~n12617;
  assign n12850 = n12849 ^ n12467;
  assign n12851 = n12850 ^ n12847;
  assign n12852 = n12848 & ~n12851;
  assign n12853 = n12852 ^ n2980;
  assign n12854 = n12853 ^ n2782;
  assign n12855 = n12471 & ~n12617;
  assign n12856 = n12855 ^ n12473;
  assign n12857 = n12856 ^ n12853;
  assign n12858 = n12854 & n12857;
  assign n12859 = n12858 ^ n2782;
  assign n12860 = n12859 ^ n2583;
  assign n12861 = n12477 & ~n12617;
  assign n12862 = n12861 ^ n12479;
  assign n12863 = n12862 ^ n12859;
  assign n12864 = n12860 & ~n12863;
  assign n12865 = n12864 ^ n2583;
  assign n12866 = n12865 ^ n2374;
  assign n12867 = n12483 & ~n12617;
  assign n12868 = n12867 ^ n12485;
  assign n12869 = n12868 ^ n12865;
  assign n12870 = n12866 & n12869;
  assign n12871 = n12870 ^ n2374;
  assign n12872 = n12871 ^ n12695;
  assign n12873 = ~n12696 & ~n12872;
  assign n12874 = n12873 ^ n2194;
  assign n12875 = n12874 ^ n12691;
  assign n12876 = ~n12692 & ~n12875;
  assign n12877 = n12876 ^ n2011;
  assign n12878 = n12877 ^ n1804;
  assign n12879 = ~n12495 & ~n12617;
  assign n12880 = n12879 ^ n12497;
  assign n12881 = n12880 ^ n12877;
  assign n12882 = n12878 & ~n12881;
  assign n12883 = n12882 ^ n1804;
  assign n12884 = n12883 ^ n1621;
  assign n12885 = n12501 & ~n12617;
  assign n12886 = n12885 ^ n12503;
  assign n12887 = n12886 ^ n12883;
  assign n12888 = n12884 & n12887;
  assign n12889 = n12888 ^ n1621;
  assign n12890 = n12889 ^ n1458;
  assign n12891 = n12507 & ~n12617;
  assign n12892 = n12891 ^ n12509;
  assign n12893 = n12892 ^ n12889;
  assign n12894 = n12890 & ~n12893;
  assign n12895 = n12894 ^ n1458;
  assign n12896 = n12895 ^ n1299;
  assign n12897 = n12513 & ~n12617;
  assign n12898 = n12897 ^ n12515;
  assign n12899 = n12898 ^ n12895;
  assign n12900 = n12896 & n12899;
  assign n12901 = n12900 ^ n1299;
  assign n12902 = n12901 ^ n1158;
  assign n12903 = n12519 & ~n12617;
  assign n12904 = n12903 ^ n12521;
  assign n12905 = n12904 ^ n12901;
  assign n12906 = n12902 & ~n12905;
  assign n12907 = n12906 ^ n1158;
  assign n12908 = n12907 ^ n1027;
  assign n12909 = n12525 & ~n12617;
  assign n12910 = n12909 ^ n12527;
  assign n12911 = n12910 ^ n12907;
  assign n12912 = n12908 & n12911;
  assign n12913 = n12912 ^ n1027;
  assign n12914 = n12913 ^ n905;
  assign n12915 = n12531 & ~n12617;
  assign n12916 = n12915 ^ n12533;
  assign n12917 = n12916 ^ n12913;
  assign n12918 = n12914 & ~n12917;
  assign n12919 = n12918 ^ n905;
  assign n12920 = n12919 ^ n803;
  assign n12921 = n12537 & ~n12617;
  assign n12922 = n12921 ^ n12539;
  assign n12923 = n12922 ^ n12919;
  assign n12924 = n12920 & n12923;
  assign n12925 = n12924 ^ n803;
  assign n12926 = n12925 ^ n707;
  assign n12927 = n12543 & ~n12617;
  assign n12928 = n12927 ^ n12545;
  assign n12929 = n12928 ^ n12925;
  assign n12930 = ~n12926 & ~n12929;
  assign n12931 = n12930 ^ n707;
  assign n12932 = n12931 ^ n608;
  assign n12933 = ~n12549 & ~n12617;
  assign n12934 = n12933 ^ n12551;
  assign n12935 = n12934 ^ n12931;
  assign n12936 = ~n12932 & ~n12935;
  assign n12937 = n12936 ^ n608;
  assign n12938 = n12937 ^ n514;
  assign n12939 = ~n12555 & ~n12617;
  assign n12940 = n12939 ^ n12557;
  assign n12941 = n12940 ^ n12937;
  assign n12942 = n12938 & ~n12941;
  assign n12943 = n12942 ^ n514;
  assign n12944 = n12943 ^ n436;
  assign n12945 = n12560 ^ n514;
  assign n12946 = ~n12617 & n12945;
  assign n12947 = n12946 ^ n12272;
  assign n12948 = n12947 ^ n12943;
  assign n12949 = n12944 & n12948;
  assign n12950 = n12949 ^ n436;
  assign n12951 = n12950 ^ n363;
  assign n12952 = ~n12561 & ~n12563;
  assign n12953 = n12952 ^ n436;
  assign n12954 = ~n12617 & n12953;
  assign n12955 = n12954 ^ n12264;
  assign n12956 = n12955 ^ n12950;
  assign n12957 = n12951 & ~n12956;
  assign n12958 = n12957 ^ n363;
  assign n12959 = n12958 ^ n300;
  assign n12960 = ~n12561 & n12564;
  assign n12961 = ~n12265 & ~n12960;
  assign n12962 = n12961 ^ n363;
  assign n12963 = ~n12617 & ~n12962;
  assign n12964 = n12963 ^ n12261;
  assign n12965 = n12964 ^ n12958;
  assign n12966 = n12959 & n12965;
  assign n12967 = n12966 ^ n300;
  assign n12968 = n12967 ^ n243;
  assign n12969 = n12961 ^ n12261;
  assign n12970 = ~n12262 & ~n12969;
  assign n12971 = n12970 ^ n363;
  assign n12972 = n12971 ^ n300;
  assign n12973 = ~n12617 & n12972;
  assign n12974 = n12973 ^ n12257;
  assign n12975 = n12974 ^ n12967;
  assign n12976 = n12968 & ~n12975;
  assign n12977 = n12976 ^ n243;
  assign n12978 = n12977 ^ n12687;
  assign n12979 = ~n12688 & n12978;
  assign n12980 = n12979 ^ n210;
  assign n12981 = n12980 ^ n12684;
  assign n12982 = ~n12685 & ~n12981;
  assign n12983 = n12982 ^ n147;
  assign n12984 = n132 & n12983;
  assign n12985 = n12579 ^ n12249;
  assign n12986 = n12682 & ~n12985;
  assign n12987 = n12986 ^ n210;
  assign n12988 = n12987 ^ n147;
  assign n12989 = ~n12617 & ~n12988;
  assign n12990 = n12989 ^ n12252;
  assign n12991 = ~n12984 & ~n12990;
  assign n12992 = ~n132 & ~n12983;
  assign n12993 = ~n12991 & ~n12992;
  assign n12994 = n12592 ^ n132;
  assign n12995 = ~n12617 & ~n12994;
  assign n12996 = n12995 ^ n12583;
  assign n12997 = ~n133 & ~n12996;
  assign n12998 = ~n12993 & ~n12997;
  assign n12999 = n12616 ^ n12591;
  assign n13000 = n12999 ^ n12591;
  assign n13001 = n12593 ^ n12591;
  assign n13002 = n13001 ^ n12591;
  assign n13003 = ~n13000 & n13002;
  assign n13004 = n13003 ^ n12591;
  assign n13005 = n12597 & ~n13004;
  assign n13006 = n13005 ^ n12591;
  assign n13007 = n133 & ~n13006;
  assign n13008 = ~n12590 & ~n12593;
  assign n13009 = ~n132 & ~n13008;
  assign n13010 = n13007 & ~n13009;
  assign n13011 = ~n12583 & n12616;
  assign n13012 = ~n12597 & n13011;
  assign n13013 = ~n13010 & ~n13012;
  assign n13014 = ~n12594 & ~n12597;
  assign n13015 = ~n12597 & ~n12616;
  assign n13016 = n12583 & ~n13015;
  assign n13017 = n13016 ^ n12592;
  assign n13018 = n13016 ^ n12597;
  assign n13019 = n13016 ^ n12994;
  assign n13020 = ~n13016 & ~n13019;
  assign n13021 = n13020 ^ n13016;
  assign n13022 = n13018 & ~n13021;
  assign n13023 = n13022 ^ n13020;
  assign n13024 = n13023 ^ n13016;
  assign n13025 = n13024 ^ n12994;
  assign n13026 = n13017 & ~n13025;
  assign n13027 = n13026 ^ n13016;
  assign n13028 = ~n13014 & ~n13027;
  assign n13029 = ~n133 & ~n13028;
  assign n13030 = n13013 & ~n13029;
  assign n13031 = ~n12998 & ~n13030;
  assign n13032 = n12681 & ~n13031;
  assign n13033 = n13032 ^ n12705;
  assign n13034 = n13033 ^ n9502;
  assign n13035 = ~n12675 & ~n13031;
  assign n13036 = n13035 ^ n12677;
  assign n13037 = n13036 ^ n9867;
  assign n13038 = n12671 ^ n10585;
  assign n13039 = ~n13031 & ~n13038;
  assign n13040 = n13039 ^ n12619;
  assign n13041 = n13040 ^ n10229;
  assign n13042 = n12635 & ~n13031;
  assign n13043 = n13042 ^ n12639;
  assign n13044 = ~n11395 & ~n13043;
  assign n13045 = n12643 & ~n13031;
  assign n13046 = n13045 ^ n12665;
  assign n13047 = ~n10956 & ~n13046;
  assign n13048 = ~n13044 & ~n13047;
  assign n13049 = x14 & n12617;
  assign n13050 = ~x12 & ~x13;
  assign n13051 = n12617 & ~n13050;
  assign n13052 = ~n13049 & ~n13051;
  assign n13053 = n13031 ^ x15;
  assign n13054 = n13052 & n13053;
  assign n13056 = ~n12617 & n13050;
  assign n13055 = ~x15 & ~n13031;
  assign n13057 = n13056 ^ n13055;
  assign n13058 = ~x14 & n13057;
  assign n13059 = n13058 ^ n13055;
  assign n13060 = ~n13054 & ~n13059;
  assign n13061 = n13060 ^ n12230;
  assign n13062 = n12624 ^ n12617;
  assign n13063 = ~n13031 & ~n13062;
  assign n13064 = n13063 ^ n12617;
  assign n13065 = n13064 ^ x16;
  assign n13066 = n13065 ^ n13060;
  assign n13067 = n13061 & n13066;
  assign n13068 = n13067 ^ n12230;
  assign n13069 = n13068 ^ n11820;
  assign n13071 = n12617 ^ n12230;
  assign n13072 = n13071 ^ n12617;
  assign n13073 = n13072 ^ n13071;
  assign n13074 = n13071 ^ n12624;
  assign n13075 = n13073 & n13074;
  assign n13076 = n13075 ^ n13071;
  assign n13077 = ~x16 & n13076;
  assign n13078 = n13077 ^ n13071;
  assign n13070 = ~x16 & ~n12617;
  assign n13079 = n13078 ^ n13070;
  assign n13080 = n12624 ^ n12230;
  assign n13081 = n13080 ^ n13078;
  assign n13082 = n13078 ^ n13031;
  assign n13083 = ~n13078 & n13082;
  assign n13084 = n13083 ^ n13078;
  assign n13085 = ~n13081 & ~n13084;
  assign n13086 = n13085 ^ n13083;
  assign n13087 = n13086 ^ n13078;
  assign n13088 = n13087 ^ n13031;
  assign n13089 = n13079 & n13088;
  assign n13090 = n13089 ^ n13070;
  assign n13091 = n13090 ^ x17;
  assign n13092 = n13091 ^ n13068;
  assign n13093 = n13069 & ~n13092;
  assign n13094 = n13093 ^ n11820;
  assign n13095 = n13048 & n13094;
  assign n13096 = n13046 ^ n10956;
  assign n13097 = n11395 & n13043;
  assign n13098 = n13097 ^ n13046;
  assign n13099 = n13096 & ~n13098;
  assign n13100 = n13099 ^ n10956;
  assign n13101 = ~n13095 & ~n13100;
  assign n13102 = n13101 ^ n10585;
  assign n13103 = n12668 ^ n10956;
  assign n13104 = ~n13031 & n13103;
  assign n13105 = n13104 ^ n12622;
  assign n13106 = n13105 ^ n13101;
  assign n13107 = n13102 & ~n13106;
  assign n13108 = n13107 ^ n10585;
  assign n13109 = n13108 ^ n13040;
  assign n13110 = n13041 & n13109;
  assign n13111 = n13110 ^ n10229;
  assign n13112 = n13111 ^ n13036;
  assign n13113 = ~n13037 & n13112;
  assign n13114 = n13113 ^ n9867;
  assign n13115 = n13114 ^ n13033;
  assign n13116 = n13034 & ~n13115;
  assign n13117 = n13116 ^ n9502;
  assign n13118 = n13117 ^ n9129;
  assign n13119 = n12983 ^ n132;
  assign n13120 = ~n13031 & n13119;
  assign n13121 = n13120 ^ n12990;
  assign n13122 = ~n133 & n13121;
  assign n13123 = n12968 & ~n13031;
  assign n13124 = n13123 ^ n12974;
  assign n13125 = ~n210 & ~n13124;
  assign n13126 = n12959 & ~n13031;
  assign n13127 = n13126 ^ n12964;
  assign n13128 = ~n243 & n13127;
  assign n13129 = ~n13125 & ~n13128;
  assign n13130 = ~n12932 & ~n13031;
  assign n13131 = n13130 ^ n12934;
  assign n13132 = n514 & ~n13131;
  assign n13133 = n12938 & ~n13031;
  assign n13134 = n13133 ^ n12940;
  assign n13135 = n436 & n13134;
  assign n13136 = ~n13132 & ~n13135;
  assign n13137 = n12884 & ~n13031;
  assign n13138 = n13137 ^ n12886;
  assign n13139 = n13138 ^ n1458;
  assign n13140 = n12878 & ~n13031;
  assign n13141 = n13140 ^ n12880;
  assign n13142 = n13141 ^ n1621;
  assign n13143 = n12874 ^ n2011;
  assign n13144 = ~n13031 & ~n13143;
  assign n13145 = n13144 ^ n12691;
  assign n13146 = n13145 ^ n1804;
  assign n13147 = n12871 ^ n2194;
  assign n13148 = ~n13031 & ~n13147;
  assign n13149 = n13148 ^ n12695;
  assign n13150 = n13149 ^ n2011;
  assign n13151 = n12770 & ~n13031;
  assign n13152 = n13151 ^ n12772;
  assign n13153 = n5625 & n13152;
  assign n13154 = n12746 & ~n13031;
  assign n13155 = n13154 ^ n12748;
  assign n13156 = ~n6802 & ~n13155;
  assign n13157 = n12740 & ~n13031;
  assign n13158 = n13157 ^ n12742;
  assign n13159 = ~n7135 & n13158;
  assign n13160 = ~n13156 & ~n13159;
  assign n13161 = n12722 & ~n13031;
  assign n13162 = n13161 ^ n12724;
  assign n13163 = n8422 & n13162;
  assign n13164 = n12727 ^ n8422;
  assign n13165 = ~n13031 & n13164;
  assign n13166 = n13165 ^ n12701;
  assign n13167 = n8083 & n13166;
  assign n13168 = ~n13163 & ~n13167;
  assign n13169 = n12709 & ~n13031;
  assign n13170 = n13169 ^ n12712;
  assign n13171 = n13170 ^ n13117;
  assign n13172 = n13118 & n13171;
  assign n13173 = n13172 ^ n9129;
  assign n13174 = n13173 ^ n8769;
  assign n13175 = n12716 & ~n13031;
  assign n13176 = n13175 ^ n12718;
  assign n13177 = n13176 ^ n13173;
  assign n13178 = n13174 & ~n13177;
  assign n13179 = n13178 ^ n8769;
  assign n13180 = n13168 & ~n13179;
  assign n13181 = n13166 ^ n8083;
  assign n13182 = ~n8422 & ~n13162;
  assign n13183 = n13182 ^ n13166;
  assign n13184 = n13181 & n13183;
  assign n13185 = n13184 ^ n8083;
  assign n13186 = ~n13180 & n13185;
  assign n13187 = n13186 ^ n7777;
  assign n13188 = n12730 ^ n8083;
  assign n13189 = ~n13031 & n13188;
  assign n13190 = n13189 ^ n12698;
  assign n13191 = n13190 ^ n13186;
  assign n13192 = n13187 & n13191;
  assign n13193 = n13192 ^ n7777;
  assign n13194 = n13193 ^ n7463;
  assign n13195 = n12734 & ~n13031;
  assign n13196 = n13195 ^ n12736;
  assign n13197 = n13196 ^ n13193;
  assign n13198 = n13194 & ~n13197;
  assign n13199 = n13198 ^ n7463;
  assign n13200 = n13160 & n13199;
  assign n13201 = n13155 ^ n6802;
  assign n13202 = n7135 & ~n13158;
  assign n13203 = n13202 ^ n13155;
  assign n13204 = n13201 & ~n13203;
  assign n13205 = n13204 ^ n6802;
  assign n13206 = ~n13200 & ~n13205;
  assign n13207 = n13206 ^ n6479;
  assign n13208 = n12752 & ~n13031;
  assign n13209 = n13208 ^ n12754;
  assign n13210 = n13209 ^ n13206;
  assign n13211 = ~n13207 & ~n13210;
  assign n13212 = n13211 ^ n6479;
  assign n13213 = n13212 ^ n6181;
  assign n13214 = n12758 & ~n13031;
  assign n13215 = n13214 ^ n12760;
  assign n13216 = n13215 ^ n13212;
  assign n13217 = n13213 & ~n13216;
  assign n13218 = n13217 ^ n6181;
  assign n13219 = n13218 ^ n5905;
  assign n13220 = n12764 & ~n13031;
  assign n13221 = n13220 ^ n12766;
  assign n13222 = n13221 ^ n13218;
  assign n13223 = n13219 & n13222;
  assign n13224 = n13223 ^ n5905;
  assign n13225 = ~n13153 & ~n13224;
  assign n13226 = ~n5625 & ~n13152;
  assign n13227 = ~n13225 & ~n13226;
  assign n13228 = n12776 & ~n13031;
  assign n13229 = n13228 ^ n12779;
  assign n13230 = n13229 ^ n5108;
  assign n13231 = n13229 ^ n5363;
  assign n13232 = n13231 ^ n5363;
  assign n13233 = n12783 & ~n13031;
  assign n13234 = n13233 ^ n12786;
  assign n13235 = n13234 ^ n5363;
  assign n13236 = ~n13232 & ~n13235;
  assign n13237 = n13236 ^ n5363;
  assign n13238 = ~n13230 & ~n13237;
  assign n13239 = n13238 ^ n5108;
  assign n13240 = n13227 & n13239;
  assign n13241 = n5363 & n13234;
  assign n13242 = ~n13226 & n13241;
  assign n13243 = ~n13225 & n13242;
  assign n13244 = n13234 ^ n5108;
  assign n13245 = n5363 & ~n13229;
  assign n13246 = n13245 ^ n13234;
  assign n13247 = n13244 & ~n13246;
  assign n13248 = n13247 ^ n5108;
  assign n13249 = ~n13243 & ~n13248;
  assign n13250 = ~n13240 & n13249;
  assign n13251 = n13250 ^ n4851;
  assign n13252 = n12790 & ~n13031;
  assign n13253 = n13252 ^ n12792;
  assign n13254 = n13253 ^ n13250;
  assign n13255 = ~n13251 & ~n13254;
  assign n13256 = n13255 ^ n4851;
  assign n13257 = n13256 ^ n4606;
  assign n13258 = n12796 & ~n13031;
  assign n13259 = n13258 ^ n12798;
  assign n13260 = n13259 ^ n13256;
  assign n13261 = n13257 & ~n13260;
  assign n13262 = n13261 ^ n4606;
  assign n13263 = n13262 ^ n4362;
  assign n13264 = n12802 & ~n13031;
  assign n13265 = n13264 ^ n12805;
  assign n13266 = n13265 ^ n13262;
  assign n13267 = n13263 & n13266;
  assign n13268 = n13267 ^ n4362;
  assign n13269 = n13268 ^ n4133;
  assign n13270 = n12809 & ~n13031;
  assign n13271 = n13270 ^ n12812;
  assign n13272 = n13271 ^ n13268;
  assign n13273 = n13269 & ~n13272;
  assign n13274 = n13273 ^ n4133;
  assign n13275 = n13274 ^ n3882;
  assign n13276 = n12816 & ~n13031;
  assign n13277 = n13276 ^ n12818;
  assign n13278 = n13277 ^ n13274;
  assign n13279 = n13275 & ~n13278;
  assign n13280 = n13279 ^ n3882;
  assign n13281 = n13280 ^ n3634;
  assign n13282 = n12822 & ~n13031;
  assign n13283 = n13282 ^ n12824;
  assign n13284 = n13283 ^ n13280;
  assign n13285 = ~n13281 & ~n13284;
  assign n13286 = n13285 ^ n3634;
  assign n13287 = n13286 ^ n3397;
  assign n13288 = ~n12828 & ~n13031;
  assign n13289 = n13288 ^ n12831;
  assign n13290 = n13289 ^ n13286;
  assign n13291 = ~n13287 & ~n13290;
  assign n13292 = n13291 ^ n3397;
  assign n13293 = n13292 ^ n3177;
  assign n13294 = ~n12835 & ~n13031;
  assign n13295 = n13294 ^ n12838;
  assign n13296 = n13295 ^ n13292;
  assign n13297 = n13293 & ~n13296;
  assign n13298 = n13297 ^ n3177;
  assign n13299 = n13298 ^ n2980;
  assign n13300 = n12842 & ~n13031;
  assign n13301 = n13300 ^ n12844;
  assign n13302 = n13301 ^ n13298;
  assign n13303 = n13299 & n13302;
  assign n13304 = n13303 ^ n2980;
  assign n13305 = n13304 ^ n2782;
  assign n13306 = n12848 & ~n13031;
  assign n13307 = n13306 ^ n12850;
  assign n13308 = n13307 ^ n13304;
  assign n13309 = n13305 & ~n13308;
  assign n13310 = n13309 ^ n2782;
  assign n13311 = n13310 ^ n2583;
  assign n13312 = n12854 & ~n13031;
  assign n13313 = n13312 ^ n12856;
  assign n13314 = n13313 ^ n13310;
  assign n13315 = n13311 & n13314;
  assign n13316 = n13315 ^ n2583;
  assign n13317 = n13316 ^ n2374;
  assign n13318 = n12860 & ~n13031;
  assign n13319 = n13318 ^ n12862;
  assign n13320 = n13319 ^ n13316;
  assign n13321 = n13317 & ~n13320;
  assign n13322 = n13321 ^ n2374;
  assign n13323 = n13322 ^ n2194;
  assign n13324 = n12866 & ~n13031;
  assign n13325 = n13324 ^ n12868;
  assign n13326 = n13325 ^ n13322;
  assign n13327 = ~n13323 & n13326;
  assign n13328 = n13327 ^ n2194;
  assign n13329 = n13328 ^ n13149;
  assign n13330 = n13150 & n13329;
  assign n13331 = n13330 ^ n2011;
  assign n13332 = n13331 ^ n13145;
  assign n13333 = ~n13146 & n13332;
  assign n13334 = n13333 ^ n1804;
  assign n13335 = n13334 ^ n13141;
  assign n13336 = n13142 & ~n13335;
  assign n13337 = n13336 ^ n1621;
  assign n13338 = n13337 ^ n13138;
  assign n13339 = ~n13139 & n13338;
  assign n13340 = n13339 ^ n1458;
  assign n13341 = n13340 ^ n1299;
  assign n13342 = n12890 & ~n13031;
  assign n13343 = n13342 ^ n12892;
  assign n13344 = n13343 ^ n13340;
  assign n13345 = n13341 & ~n13344;
  assign n13346 = n13345 ^ n1299;
  assign n13347 = n13346 ^ n1158;
  assign n13348 = n12896 & ~n13031;
  assign n13349 = n13348 ^ n12898;
  assign n13350 = n13349 ^ n13346;
  assign n13351 = n13347 & n13350;
  assign n13352 = n13351 ^ n1158;
  assign n13353 = n13352 ^ n1027;
  assign n13354 = n12902 & ~n13031;
  assign n13355 = n13354 ^ n12904;
  assign n13356 = n13355 ^ n13352;
  assign n13357 = n13353 & ~n13356;
  assign n13358 = n13357 ^ n1027;
  assign n13359 = n13358 ^ n905;
  assign n13360 = n12908 & ~n13031;
  assign n13361 = n13360 ^ n12910;
  assign n13362 = n13361 ^ n13358;
  assign n13363 = n13359 & n13362;
  assign n13364 = n13363 ^ n905;
  assign n13365 = n13364 ^ n803;
  assign n13366 = n12914 & ~n13031;
  assign n13367 = n13366 ^ n12916;
  assign n13368 = n13367 ^ n13364;
  assign n13369 = n13365 & ~n13368;
  assign n13370 = n13369 ^ n803;
  assign n13371 = n13370 ^ n707;
  assign n13372 = n12920 & ~n13031;
  assign n13373 = n13372 ^ n12922;
  assign n13374 = n13373 ^ n13370;
  assign n13375 = ~n13371 & n13374;
  assign n13376 = n13375 ^ n707;
  assign n13377 = n13376 ^ n608;
  assign n13378 = ~n12926 & ~n13031;
  assign n13379 = n13378 ^ n12928;
  assign n13380 = n13379 ^ n13376;
  assign n13381 = ~n13377 & n13380;
  assign n13382 = n13381 ^ n608;
  assign n13383 = n13136 & ~n13382;
  assign n13384 = n13134 ^ n436;
  assign n13385 = ~n514 & n13131;
  assign n13386 = n13385 ^ n13134;
  assign n13387 = n13384 & n13386;
  assign n13388 = n13387 ^ n436;
  assign n13389 = ~n13383 & n13388;
  assign n13390 = n13389 ^ n363;
  assign n13391 = n12944 & ~n13031;
  assign n13392 = n13391 ^ n12947;
  assign n13393 = n13392 ^ n13389;
  assign n13394 = n13390 & n13393;
  assign n13395 = n13394 ^ n363;
  assign n13396 = n13395 ^ n300;
  assign n13397 = n12951 & ~n13031;
  assign n13398 = n13397 ^ n12955;
  assign n13399 = n13398 ^ n13395;
  assign n13400 = n13396 & ~n13399;
  assign n13401 = n13400 ^ n300;
  assign n13402 = n13129 & n13401;
  assign n13403 = n13124 ^ n210;
  assign n13404 = n243 & ~n13127;
  assign n13405 = n13404 ^ n13124;
  assign n13406 = n13403 & ~n13405;
  assign n13407 = n13406 ^ n210;
  assign n13408 = ~n13402 & ~n13407;
  assign n13409 = n13408 ^ n147;
  assign n13410 = n12977 ^ n210;
  assign n13411 = ~n13031 & n13410;
  assign n13412 = n13411 ^ n12687;
  assign n13413 = n13412 ^ n13408;
  assign n13414 = n13409 & ~n13413;
  assign n13415 = n13414 ^ n147;
  assign n13416 = n13415 ^ n132;
  assign n13417 = n12980 ^ n147;
  assign n13418 = ~n13031 & ~n13417;
  assign n13419 = n13418 ^ n12684;
  assign n13420 = n13419 ^ n13415;
  assign n13421 = n13416 & n13420;
  assign n13422 = n13421 ^ n132;
  assign n13423 = ~n13122 & ~n13422;
  assign n13424 = ~n133 & ~n12993;
  assign n13425 = n1292 & n13030;
  assign n13426 = n12990 & n13425;
  assign n13427 = n12983 & n13426;
  assign n13428 = n12996 & ~n13427;
  assign n13429 = ~n13424 & n13428;
  assign n13434 = n12997 & n13030;
  assign n13430 = ~n12992 & n13030;
  assign n13431 = n12990 & ~n13430;
  assign n13432 = n133 & ~n12996;
  assign n13433 = ~n13431 & n13432;
  assign n13435 = n13434 ^ n13433;
  assign n13436 = n12992 ^ n12991;
  assign n13437 = n13436 ^ n12991;
  assign n13438 = n13434 ^ n12991;
  assign n13439 = n13437 & n13438;
  assign n13440 = n13439 ^ n12991;
  assign n13441 = n13435 & n13440;
  assign n13442 = n13441 ^ n13433;
  assign n13443 = ~n13429 & ~n13442;
  assign n13444 = ~n13423 & n13443;
  assign n13445 = n13118 & ~n13444;
  assign n13446 = n13445 ^ n13170;
  assign n13447 = n13446 ^ n8769;
  assign n13448 = n13114 ^ n9502;
  assign n13449 = ~n13444 & n13448;
  assign n13450 = n13449 ^ n13033;
  assign n13451 = n13450 ^ n9129;
  assign n13452 = ~x10 & ~x11;
  assign n13453 = ~x12 & n13452;
  assign n13454 = n13031 & ~n13453;
  assign n13455 = n13444 ^ x13;
  assign n13456 = ~n13454 & n13455;
  assign n13458 = ~n13031 & n13452;
  assign n13457 = ~x13 & ~n13444;
  assign n13459 = n13458 ^ n13457;
  assign n13460 = ~x12 & n13459;
  assign n13461 = n13460 ^ n13457;
  assign n13462 = ~n13456 & ~n13461;
  assign n13463 = n13462 ^ n12617;
  assign n13464 = n13050 ^ n13031;
  assign n13465 = ~n13444 & ~n13464;
  assign n13466 = n13465 ^ n13031;
  assign n13467 = n13466 ^ x14;
  assign n13468 = n13467 ^ n13462;
  assign n13469 = n13463 & n13468;
  assign n13470 = n13469 ^ n12617;
  assign n13471 = n13470 ^ n12230;
  assign n13473 = ~x14 & n13050;
  assign n13474 = n13473 ^ n12617;
  assign n13475 = n13474 ^ n13049;
  assign n13476 = n13031 & ~n13475;
  assign n13477 = n13476 ^ n13049;
  assign n13472 = ~x14 & ~n13031;
  assign n13478 = n13477 ^ n13472;
  assign n13479 = n13050 ^ n12617;
  assign n13480 = n13479 ^ n13477;
  assign n13481 = n13477 ^ n13444;
  assign n13482 = ~n13477 & n13481;
  assign n13483 = n13482 ^ n13477;
  assign n13484 = ~n13480 & ~n13483;
  assign n13485 = n13484 ^ n13482;
  assign n13486 = n13485 ^ n13477;
  assign n13487 = n13486 ^ n13444;
  assign n13488 = n13478 & n13487;
  assign n13489 = n13488 ^ n13472;
  assign n13490 = n13489 ^ x15;
  assign n13491 = n13490 ^ n13470;
  assign n13492 = n13471 & ~n13491;
  assign n13493 = n13492 ^ n12230;
  assign n13494 = n13493 ^ n11820;
  assign n13495 = n13061 & ~n13444;
  assign n13496 = n13495 ^ n13065;
  assign n13497 = n13496 ^ n13493;
  assign n13498 = n13494 & n13497;
  assign n13499 = n13498 ^ n11820;
  assign n13500 = n13499 ^ n11395;
  assign n13501 = n13069 & ~n13444;
  assign n13502 = n13501 ^ n13091;
  assign n13503 = n13502 ^ n13499;
  assign n13504 = n13500 & ~n13503;
  assign n13505 = n13504 ^ n11395;
  assign n13506 = n13505 ^ n10956;
  assign n13507 = n13094 ^ n11395;
  assign n13508 = ~n13444 & n13507;
  assign n13509 = n13508 ^ n13043;
  assign n13510 = n13509 ^ n13505;
  assign n13511 = n13506 & ~n13510;
  assign n13512 = n13511 ^ n10956;
  assign n13513 = n13512 ^ n10585;
  assign n13514 = n13094 ^ n13043;
  assign n13515 = n13507 & ~n13514;
  assign n13516 = n13515 ^ n11395;
  assign n13517 = n13516 ^ n10956;
  assign n13518 = ~n13444 & n13517;
  assign n13519 = n13518 ^ n13046;
  assign n13520 = n13519 ^ n13512;
  assign n13521 = ~n13513 & ~n13520;
  assign n13522 = n13521 ^ n10585;
  assign n13523 = n13522 ^ n10229;
  assign n13524 = n13102 & ~n13444;
  assign n13525 = n13524 ^ n13105;
  assign n13526 = n13525 ^ n13522;
  assign n13527 = ~n13523 & ~n13526;
  assign n13528 = n13527 ^ n10229;
  assign n13529 = n13528 ^ n9867;
  assign n13530 = n13108 ^ n10229;
  assign n13531 = ~n13444 & ~n13530;
  assign n13532 = n13531 ^ n13040;
  assign n13533 = n13532 ^ n13528;
  assign n13534 = n13529 & ~n13533;
  assign n13535 = n13534 ^ n9867;
  assign n13536 = n13535 ^ n9502;
  assign n13537 = n13111 ^ n9867;
  assign n13538 = ~n13444 & n13537;
  assign n13539 = n13538 ^ n13036;
  assign n13540 = n13539 ^ n13535;
  assign n13541 = n13536 & n13540;
  assign n13542 = n13541 ^ n9502;
  assign n13543 = n13542 ^ n13450;
  assign n13544 = n13451 & ~n13543;
  assign n13545 = n13544 ^ n9129;
  assign n13546 = n13545 ^ n13446;
  assign n13547 = ~n13447 & n13546;
  assign n13548 = n13547 ^ n8769;
  assign n13549 = n13548 ^ n8422;
  assign n13550 = n13174 & ~n13444;
  assign n13551 = n13550 ^ n13176;
  assign n13552 = n13551 ^ n13548;
  assign n13553 = n13549 & ~n13552;
  assign n13554 = n13553 ^ n8422;
  assign n13555 = n13554 ^ n8083;
  assign n13556 = n13422 ^ n133;
  assign n13557 = n13556 ^ n13121;
  assign n13558 = n13443 & ~n13556;
  assign n13559 = n13557 & n13558;
  assign n13560 = n13559 ^ n13557;
  assign n13561 = n13337 ^ n1458;
  assign n13562 = ~n13444 & n13561;
  assign n13563 = n13562 ^ n13138;
  assign n13564 = n13563 ^ n1299;
  assign n13565 = n13334 ^ n1621;
  assign n13566 = ~n13444 & n13565;
  assign n13567 = n13566 ^ n13141;
  assign n13568 = n13567 ^ n1458;
  assign n13569 = n2011 & ~n2194;
  assign n13570 = n13317 & ~n13444;
  assign n13571 = n13570 ^ n13319;
  assign n13572 = ~n13569 & ~n13571;
  assign n13573 = n13269 & ~n13444;
  assign n13574 = n13573 ^ n13271;
  assign n13575 = n13574 ^ n3882;
  assign n13576 = n13263 & ~n13444;
  assign n13577 = n13576 ^ n13265;
  assign n13578 = n13577 ^ n4133;
  assign n13579 = n13224 ^ n5625;
  assign n13580 = ~n13444 & n13579;
  assign n13581 = n13580 ^ n13152;
  assign n13582 = n13581 ^ n5363;
  assign n13583 = n13219 & ~n13444;
  assign n13584 = n13583 ^ n13221;
  assign n13585 = n13584 ^ n5625;
  assign n13586 = n13179 ^ n8422;
  assign n13587 = ~n13444 & n13586;
  assign n13588 = n13587 ^ n13162;
  assign n13589 = n13588 ^ n13554;
  assign n13590 = n13555 & ~n13589;
  assign n13591 = n13590 ^ n8083;
  assign n13592 = n13591 ^ n7777;
  assign n13593 = n13179 ^ n13162;
  assign n13594 = n13586 & ~n13593;
  assign n13595 = n13594 ^ n8422;
  assign n13596 = n13595 ^ n8083;
  assign n13597 = ~n13444 & n13596;
  assign n13598 = n13597 ^ n13166;
  assign n13599 = n13598 ^ n13591;
  assign n13600 = n13592 & ~n13599;
  assign n13601 = n13600 ^ n7777;
  assign n13602 = n13601 ^ n7463;
  assign n13603 = n13187 & ~n13444;
  assign n13604 = n13603 ^ n13190;
  assign n13605 = n13604 ^ n13601;
  assign n13606 = n13602 & n13605;
  assign n13607 = n13606 ^ n7463;
  assign n13608 = n13607 ^ n7135;
  assign n13609 = n13194 & ~n13444;
  assign n13610 = n13609 ^ n13196;
  assign n13611 = n13610 ^ n13607;
  assign n13612 = n13608 & ~n13611;
  assign n13613 = n13612 ^ n7135;
  assign n13614 = n13613 ^ n6802;
  assign n13615 = n13199 ^ n7135;
  assign n13616 = ~n13444 & n13615;
  assign n13617 = n13616 ^ n13158;
  assign n13618 = n13617 ^ n13613;
  assign n13619 = n13614 & n13618;
  assign n13620 = n13619 ^ n6802;
  assign n13621 = n13620 ^ n6479;
  assign n13622 = n13199 ^ n13158;
  assign n13623 = n13615 & n13622;
  assign n13624 = n13623 ^ n7135;
  assign n13625 = n13624 ^ n6802;
  assign n13626 = ~n13444 & n13625;
  assign n13627 = n13626 ^ n13155;
  assign n13628 = n13627 ^ n13620;
  assign n13629 = n13621 & ~n13628;
  assign n13630 = n13629 ^ n6479;
  assign n13631 = n13630 ^ n6181;
  assign n13632 = ~n13207 & ~n13444;
  assign n13633 = n13632 ^ n13209;
  assign n13634 = n13633 ^ n13630;
  assign n13635 = n13631 & n13634;
  assign n13636 = n13635 ^ n6181;
  assign n13637 = n13636 ^ n5905;
  assign n13638 = n13213 & ~n13444;
  assign n13639 = n13638 ^ n13215;
  assign n13640 = n13639 ^ n13636;
  assign n13641 = n13637 & ~n13640;
  assign n13642 = n13641 ^ n5905;
  assign n13643 = n13642 ^ n13584;
  assign n13644 = ~n13585 & n13643;
  assign n13645 = n13644 ^ n5625;
  assign n13646 = n13645 ^ n13581;
  assign n13647 = n13582 & ~n13646;
  assign n13648 = n13647 ^ n5363;
  assign n13649 = n13648 ^ n5108;
  assign n13650 = n13227 ^ n5363;
  assign n13651 = ~n13444 & n13650;
  assign n13652 = n13651 ^ n13229;
  assign n13653 = n13652 ^ n13648;
  assign n13654 = n13649 & n13653;
  assign n13655 = n13654 ^ n5108;
  assign n13656 = n13655 ^ n4851;
  assign n13657 = n13229 ^ n13227;
  assign n13658 = n13650 & n13657;
  assign n13659 = n13658 ^ n5363;
  assign n13660 = n13659 ^ n5108;
  assign n13661 = ~n13444 & n13660;
  assign n13662 = n13661 ^ n13234;
  assign n13663 = n13662 ^ n13655;
  assign n13664 = n13656 & ~n13663;
  assign n13665 = n13664 ^ n4851;
  assign n13666 = n13665 ^ n4606;
  assign n13667 = ~n13251 & ~n13444;
  assign n13668 = n13667 ^ n13253;
  assign n13669 = n13668 ^ n13665;
  assign n13670 = n13666 & n13669;
  assign n13671 = n13670 ^ n4606;
  assign n13672 = n13671 ^ n4362;
  assign n13673 = n13257 & ~n13444;
  assign n13674 = n13673 ^ n13259;
  assign n13675 = n13674 ^ n13671;
  assign n13676 = n13672 & ~n13675;
  assign n13677 = n13676 ^ n4362;
  assign n13678 = n13677 ^ n13577;
  assign n13679 = ~n13578 & n13678;
  assign n13680 = n13679 ^ n4133;
  assign n13681 = n13680 ^ n13574;
  assign n13682 = n13575 & ~n13681;
  assign n13683 = n13682 ^ n3882;
  assign n13684 = n13683 ^ n3634;
  assign n13685 = n13275 & ~n13444;
  assign n13686 = n13685 ^ n13277;
  assign n13687 = n13686 ^ n13683;
  assign n13688 = ~n13684 & ~n13687;
  assign n13689 = n13688 ^ n3634;
  assign n13690 = n13689 ^ n3397;
  assign n13691 = ~n13281 & ~n13444;
  assign n13692 = n13691 ^ n13283;
  assign n13693 = n13692 ^ n13689;
  assign n13694 = ~n13690 & n13693;
  assign n13695 = n13694 ^ n3397;
  assign n13696 = n13695 ^ n3177;
  assign n13697 = ~n13287 & ~n13444;
  assign n13698 = n13697 ^ n13289;
  assign n13699 = n13698 ^ n13695;
  assign n13700 = n13696 & n13699;
  assign n13701 = n13700 ^ n3177;
  assign n13702 = n13701 ^ n2980;
  assign n13703 = n13293 & ~n13444;
  assign n13704 = n13703 ^ n13295;
  assign n13705 = n13704 ^ n13701;
  assign n13706 = n13702 & ~n13705;
  assign n13707 = n13706 ^ n2980;
  assign n13708 = n13707 ^ n2782;
  assign n13709 = n13299 & ~n13444;
  assign n13710 = n13709 ^ n13301;
  assign n13711 = n13710 ^ n13707;
  assign n13712 = n13708 & n13711;
  assign n13713 = n13712 ^ n2782;
  assign n13714 = n13713 ^ n2583;
  assign n13715 = n13305 & ~n13444;
  assign n13716 = n13715 ^ n13307;
  assign n13717 = n13716 ^ n13713;
  assign n13718 = n13714 & ~n13717;
  assign n13719 = n13718 ^ n2583;
  assign n13720 = n13719 ^ n2374;
  assign n13721 = n13311 & ~n13444;
  assign n13722 = n13721 ^ n13313;
  assign n13723 = n13722 ^ n13719;
  assign n13724 = n13720 & n13723;
  assign n13725 = n13724 ^ n2374;
  assign n13726 = ~n13572 & n13725;
  assign n13727 = ~n13323 & ~n13444;
  assign n13728 = n13727 ^ n13325;
  assign n13729 = n2011 & ~n13728;
  assign n13730 = ~n2194 & n13571;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = ~n13726 & n13731;
  assign n13733 = n13732 ^ n13728;
  assign n13734 = ~n2194 & n13725;
  assign n13735 = n13734 ^ n13732;
  assign n13736 = n13735 ^ n13734;
  assign n13737 = n13734 ^ n2011;
  assign n13738 = ~n13736 & ~n13737;
  assign n13739 = n13738 ^ n13734;
  assign n13740 = n13733 & ~n13739;
  assign n13741 = n13740 ^ n13728;
  assign n13742 = n13741 ^ n1804;
  assign n13743 = n13328 ^ n2011;
  assign n13744 = ~n13444 & ~n13743;
  assign n13745 = n13744 ^ n13149;
  assign n13746 = n13745 ^ n13741;
  assign n13747 = ~n13742 & n13746;
  assign n13748 = n13747 ^ n1804;
  assign n13749 = n13748 ^ n1621;
  assign n13750 = n13331 ^ n1804;
  assign n13751 = ~n13444 & n13750;
  assign n13752 = n13751 ^ n13145;
  assign n13753 = n13752 ^ n13748;
  assign n13754 = n13749 & n13753;
  assign n13755 = n13754 ^ n1621;
  assign n13756 = n13755 ^ n13567;
  assign n13757 = n13568 & ~n13756;
  assign n13758 = n13757 ^ n1458;
  assign n13759 = n13758 ^ n13563;
  assign n13760 = ~n13564 & n13759;
  assign n13761 = n13760 ^ n1299;
  assign n13762 = n13761 ^ n1158;
  assign n13763 = n13341 & ~n13444;
  assign n13764 = n13763 ^ n13343;
  assign n13765 = n13764 ^ n13761;
  assign n13766 = n13762 & ~n13765;
  assign n13767 = n13766 ^ n1158;
  assign n13768 = n13767 ^ n1027;
  assign n13769 = n13347 & ~n13444;
  assign n13770 = n13769 ^ n13349;
  assign n13771 = n13770 ^ n13767;
  assign n13772 = n13768 & n13771;
  assign n13773 = n13772 ^ n1027;
  assign n13774 = n13773 ^ n905;
  assign n13775 = n13353 & ~n13444;
  assign n13776 = n13775 ^ n13355;
  assign n13777 = n13776 ^ n13773;
  assign n13778 = n13774 & ~n13777;
  assign n13779 = n13778 ^ n905;
  assign n13780 = n13779 ^ n803;
  assign n13781 = n13359 & ~n13444;
  assign n13782 = n13781 ^ n13361;
  assign n13783 = n13782 ^ n13779;
  assign n13784 = n13780 & n13783;
  assign n13785 = n13784 ^ n803;
  assign n13786 = n13785 ^ n707;
  assign n13787 = n13365 & ~n13444;
  assign n13788 = n13787 ^ n13367;
  assign n13789 = n13788 ^ n13785;
  assign n13790 = ~n13786 & ~n13789;
  assign n13791 = n13790 ^ n707;
  assign n13792 = n13791 ^ n608;
  assign n13793 = ~n13371 & ~n13444;
  assign n13794 = n13793 ^ n13373;
  assign n13795 = n13794 ^ n13791;
  assign n13796 = ~n13792 & ~n13795;
  assign n13797 = n13796 ^ n608;
  assign n13798 = n13797 ^ n514;
  assign n13799 = ~n13377 & ~n13444;
  assign n13800 = n13799 ^ n13379;
  assign n13801 = n13800 ^ n13797;
  assign n13802 = n13798 & ~n13801;
  assign n13803 = n13802 ^ n514;
  assign n13804 = n13803 ^ n436;
  assign n13805 = n13382 ^ n514;
  assign n13806 = ~n13444 & n13805;
  assign n13807 = n13806 ^ n13131;
  assign n13808 = n13807 ^ n13803;
  assign n13809 = n13804 & n13808;
  assign n13810 = n13809 ^ n436;
  assign n13811 = n13810 ^ n363;
  assign n13812 = n13382 ^ n13131;
  assign n13813 = n13805 & n13812;
  assign n13814 = n13813 ^ n514;
  assign n13815 = n13814 ^ n436;
  assign n13816 = ~n13444 & n13815;
  assign n13817 = n13816 ^ n13134;
  assign n13818 = n13817 ^ n13810;
  assign n13819 = n13811 & ~n13818;
  assign n13820 = n13819 ^ n363;
  assign n13821 = n13820 ^ n300;
  assign n13822 = n13390 & ~n13444;
  assign n13823 = n13822 ^ n13392;
  assign n13824 = n13823 ^ n13820;
  assign n13825 = n13821 & n13824;
  assign n13826 = n13825 ^ n300;
  assign n13827 = n13826 ^ n243;
  assign n13828 = n13396 & ~n13444;
  assign n13829 = n13828 ^ n13398;
  assign n13830 = n13829 ^ n13826;
  assign n13831 = n13827 & ~n13830;
  assign n13832 = n13831 ^ n243;
  assign n13833 = n13832 ^ n210;
  assign n13834 = n13401 ^ n243;
  assign n13835 = ~n13444 & n13834;
  assign n13836 = n13835 ^ n13127;
  assign n13837 = n13836 ^ n13832;
  assign n13838 = n13833 & n13837;
  assign n13839 = n13838 ^ n210;
  assign n13840 = n13839 ^ n147;
  assign n13841 = n13401 ^ n13127;
  assign n13842 = n13834 & n13841;
  assign n13843 = n13842 ^ n243;
  assign n13844 = n13843 ^ n210;
  assign n13845 = ~n13444 & n13844;
  assign n13846 = n13845 ^ n13124;
  assign n13847 = n13846 ^ n13839;
  assign n13848 = ~n13840 & ~n13847;
  assign n13849 = n13848 ^ n147;
  assign n13850 = n13849 ^ n132;
  assign n13851 = n13409 & ~n13444;
  assign n13852 = n13851 ^ n13412;
  assign n13853 = n13852 ^ n13849;
  assign n13854 = n13850 & ~n13853;
  assign n13855 = n13854 ^ n132;
  assign n13856 = n13855 ^ n133;
  assign n13857 = n13416 & ~n13444;
  assign n13858 = n13857 ^ n13419;
  assign n13859 = n13858 ^ n13855;
  assign n13860 = ~n13856 & ~n13859;
  assign n13861 = n13860 ^ n13855;
  assign n13862 = ~n13560 & n13861;
  assign n13863 = n13555 & ~n13862;
  assign n13864 = n13863 ^ n13588;
  assign n13865 = ~n7777 & ~n13864;
  assign n13866 = n13549 & ~n13862;
  assign n13867 = n13866 ^ n13551;
  assign n13868 = ~n8083 & ~n13867;
  assign n13869 = ~n13865 & ~n13868;
  assign n13870 = ~x8 & ~x9;
  assign n13871 = ~x10 & n13870;
  assign n13872 = n13444 & ~n13871;
  assign n13873 = n13862 ^ x11;
  assign n13874 = ~n13872 & n13873;
  assign n13876 = ~n13444 & n13870;
  assign n13875 = ~x11 & ~n13862;
  assign n13877 = n13876 ^ n13875;
  assign n13878 = ~x10 & n13877;
  assign n13879 = n13878 ^ n13875;
  assign n13880 = ~n13874 & ~n13879;
  assign n13881 = n13880 ^ n13031;
  assign n13882 = n13452 ^ n13444;
  assign n13883 = ~n13862 & ~n13882;
  assign n13884 = n13883 ^ n13444;
  assign n13885 = n13884 ^ x12;
  assign n13886 = n13885 ^ n13880;
  assign n13887 = n13881 & n13886;
  assign n13888 = n13887 ^ n13031;
  assign n13889 = n13888 ^ n12617;
  assign n13891 = n13453 ^ n13031;
  assign n13892 = n13891 ^ x12;
  assign n13893 = n13892 ^ n13891;
  assign n13894 = n13891 ^ n13453;
  assign n13895 = n13893 & n13894;
  assign n13896 = n13895 ^ n13891;
  assign n13897 = ~n13444 & ~n13896;
  assign n13898 = n13897 ^ n13891;
  assign n13890 = ~x12 & ~n13444;
  assign n13899 = n13898 ^ n13890;
  assign n13900 = n13452 ^ n13031;
  assign n13901 = n13900 ^ n13898;
  assign n13902 = n13898 ^ n13862;
  assign n13903 = n13898 & ~n13902;
  assign n13904 = n13903 ^ n13898;
  assign n13905 = n13901 & n13904;
  assign n13906 = n13905 ^ n13903;
  assign n13907 = n13906 ^ n13898;
  assign n13908 = n13907 ^ n13862;
  assign n13909 = ~n13899 & ~n13908;
  assign n13910 = n13909 ^ n13890;
  assign n13911 = n13910 ^ x13;
  assign n13912 = n13911 ^ n13888;
  assign n13913 = n13889 & ~n13912;
  assign n13914 = n13913 ^ n12617;
  assign n13915 = n13914 ^ n12230;
  assign n13916 = n13463 & ~n13862;
  assign n13917 = n13916 ^ n13467;
  assign n13918 = n13917 ^ n13914;
  assign n13919 = n13915 & n13918;
  assign n13920 = n13919 ^ n12230;
  assign n13921 = n13920 ^ n11820;
  assign n13922 = n13471 & ~n13862;
  assign n13923 = n13922 ^ n13490;
  assign n13924 = n13923 ^ n13920;
  assign n13925 = n13921 & ~n13924;
  assign n13926 = n13925 ^ n11820;
  assign n13927 = n13926 ^ n11395;
  assign n13928 = n13494 & ~n13862;
  assign n13929 = n13928 ^ n13496;
  assign n13930 = n13929 ^ n13926;
  assign n13931 = n13927 & n13930;
  assign n13932 = n13931 ^ n11395;
  assign n13933 = n13932 ^ n10956;
  assign n13934 = n13500 & ~n13862;
  assign n13935 = n13934 ^ n13502;
  assign n13936 = n13935 ^ n13932;
  assign n13937 = n13933 & ~n13936;
  assign n13938 = n13937 ^ n10956;
  assign n13939 = n13938 ^ n10585;
  assign n13940 = n13506 & ~n13862;
  assign n13941 = n13940 ^ n13509;
  assign n13942 = n13941 ^ n13938;
  assign n13943 = ~n13939 & ~n13942;
  assign n13944 = n13943 ^ n10585;
  assign n13945 = n13944 ^ n10229;
  assign n13946 = ~n13513 & ~n13862;
  assign n13947 = n13946 ^ n13519;
  assign n13948 = n13947 ^ n13944;
  assign n13949 = ~n13945 & n13948;
  assign n13950 = n13949 ^ n10229;
  assign n13951 = n13950 ^ n9867;
  assign n13952 = ~n13523 & ~n13862;
  assign n13953 = n13952 ^ n13525;
  assign n13954 = n13953 ^ n13950;
  assign n13955 = n13951 & n13954;
  assign n13956 = n13955 ^ n9867;
  assign n13957 = n13956 ^ n9502;
  assign n13958 = n13529 & ~n13862;
  assign n13959 = n13958 ^ n13532;
  assign n13960 = n13959 ^ n13956;
  assign n13961 = n13957 & ~n13960;
  assign n13962 = n13961 ^ n9502;
  assign n13963 = n13962 ^ n9129;
  assign n13964 = n13536 & ~n13862;
  assign n13965 = n13964 ^ n13539;
  assign n13966 = n13965 ^ n13962;
  assign n13967 = n13963 & n13966;
  assign n13968 = n13967 ^ n9129;
  assign n13969 = n13968 ^ n8769;
  assign n13970 = n13542 ^ n9129;
  assign n13971 = ~n13862 & n13970;
  assign n13972 = n13971 ^ n13450;
  assign n13973 = n13972 ^ n13968;
  assign n13974 = n13969 & ~n13973;
  assign n13975 = n13974 ^ n8769;
  assign n13976 = n13975 ^ n8422;
  assign n13977 = n13545 ^ n8769;
  assign n13978 = ~n13862 & n13977;
  assign n13979 = n13978 ^ n13446;
  assign n13980 = n13979 ^ n13975;
  assign n13981 = n13976 & n13980;
  assign n13982 = n13981 ^ n8422;
  assign n13983 = n13869 & n13982;
  assign n13984 = n13864 ^ n7777;
  assign n13985 = n8083 & n13867;
  assign n13986 = n13985 ^ n13864;
  assign n13987 = n13984 & ~n13986;
  assign n13988 = n13987 ^ n7777;
  assign n13989 = ~n13983 & ~n13988;
  assign n13990 = n13989 ^ n7463;
  assign n13991 = n13592 & ~n13862;
  assign n13992 = n13991 ^ n13598;
  assign n13993 = n13992 ^ n13989;
  assign n13994 = ~n13990 & n13993;
  assign n13995 = n13994 ^ n7463;
  assign n13996 = n13995 ^ n7135;
  assign n13997 = n13602 & ~n13862;
  assign n13998 = n13997 ^ n13604;
  assign n13999 = n13998 ^ n13995;
  assign n14000 = n13996 & n13999;
  assign n14001 = n14000 ^ n7135;
  assign n14002 = n14001 ^ n6802;
  assign n14003 = n13608 & ~n13862;
  assign n14004 = n14003 ^ n13610;
  assign n14005 = n14004 ^ n14001;
  assign n14006 = n14002 & ~n14005;
  assign n14007 = n14006 ^ n6802;
  assign n14008 = n14007 ^ n6479;
  assign n14009 = n13858 ^ n13856;
  assign n14010 = ~n13560 & ~n13856;
  assign n14011 = ~n14009 & n14010;
  assign n14012 = n14011 ^ n14009;
  assign n14015 = n13827 & ~n13862;
  assign n14016 = n14015 ^ n13829;
  assign n14017 = n14016 ^ n210;
  assign n14018 = n13821 & ~n13862;
  assign n14019 = n14018 ^ n13823;
  assign n14020 = n14019 ^ n243;
  assign n14021 = ~n13690 & ~n13862;
  assign n14022 = n14021 ^ n13692;
  assign n14023 = n13642 ^ n5625;
  assign n14024 = ~n13862 & n14023;
  assign n14025 = n14024 ^ n13584;
  assign n14026 = ~n5363 & n14025;
  assign n14027 = n13614 & ~n13862;
  assign n14028 = n14027 ^ n13617;
  assign n14029 = n14028 ^ n14007;
  assign n14030 = n14008 & n14029;
  assign n14031 = n14030 ^ n6479;
  assign n14032 = n14031 ^ n6181;
  assign n14033 = n13621 & ~n13862;
  assign n14034 = n14033 ^ n13627;
  assign n14035 = n14034 ^ n14031;
  assign n14036 = n14032 & ~n14035;
  assign n14037 = n14036 ^ n6181;
  assign n14038 = n14037 ^ n5905;
  assign n14039 = n13631 & ~n13862;
  assign n14040 = n14039 ^ n13633;
  assign n14041 = n14040 ^ n14037;
  assign n14042 = n14038 & n14041;
  assign n14043 = n14042 ^ n5905;
  assign n14044 = n14043 ^ n5625;
  assign n14045 = n13637 & ~n13862;
  assign n14046 = n14045 ^ n13639;
  assign n14047 = n14046 ^ n14043;
  assign n14048 = n14044 & ~n14047;
  assign n14049 = n14048 ^ n5625;
  assign n14050 = ~n14026 & n14049;
  assign n14051 = n5108 & n5363;
  assign n14052 = n13645 ^ n5363;
  assign n14053 = ~n13862 & n14052;
  assign n14054 = n14053 ^ n13581;
  assign n14055 = ~n14051 & ~n14054;
  assign n14056 = n14050 & ~n14055;
  assign n14057 = n5108 & ~n14025;
  assign n14058 = n14049 & n14057;
  assign n14059 = n14054 ^ n5108;
  assign n14060 = n5363 & ~n14025;
  assign n14061 = n14060 ^ n14054;
  assign n14062 = n14059 & ~n14061;
  assign n14063 = n14062 ^ n5108;
  assign n14064 = ~n14058 & ~n14063;
  assign n14065 = ~n14056 & n14064;
  assign n14066 = n14065 ^ n4851;
  assign n14067 = n13649 & ~n13862;
  assign n14068 = n14067 ^ n13652;
  assign n14069 = n14068 ^ n14065;
  assign n14070 = ~n14066 & ~n14069;
  assign n14071 = n14070 ^ n4851;
  assign n14072 = n14071 ^ n4606;
  assign n14073 = n13656 & ~n13862;
  assign n14074 = n14073 ^ n13662;
  assign n14075 = n14074 ^ n14071;
  assign n14076 = n14072 & ~n14075;
  assign n14077 = n14076 ^ n4606;
  assign n14078 = n14077 ^ n4362;
  assign n14079 = n13666 & ~n13862;
  assign n14080 = n14079 ^ n13668;
  assign n14081 = n14080 ^ n14077;
  assign n14082 = n14078 & n14081;
  assign n14083 = n14082 ^ n4362;
  assign n14084 = n14083 ^ n4133;
  assign n14085 = n13672 & ~n13862;
  assign n14086 = n14085 ^ n13674;
  assign n14087 = n14086 ^ n14083;
  assign n14088 = n14084 & ~n14087;
  assign n14089 = n14088 ^ n4133;
  assign n14090 = n14089 ^ n3882;
  assign n14091 = n13677 ^ n4133;
  assign n14092 = ~n13862 & n14091;
  assign n14093 = n14092 ^ n13577;
  assign n14094 = n14093 ^ n14089;
  assign n14095 = n14090 & n14094;
  assign n14096 = n14095 ^ n3882;
  assign n14097 = n14096 ^ n3634;
  assign n14098 = n13680 ^ n3882;
  assign n14099 = ~n13862 & n14098;
  assign n14100 = n14099 ^ n13574;
  assign n14101 = n14100 ^ n14096;
  assign n14102 = ~n14097 & ~n14101;
  assign n14103 = n14102 ^ n3634;
  assign n14104 = n14103 ^ n3397;
  assign n14105 = ~n13684 & ~n13862;
  assign n14106 = n14105 ^ n13686;
  assign n14107 = n14106 ^ n14103;
  assign n14108 = ~n14104 & n14107;
  assign n14109 = n14108 ^ n3397;
  assign n14110 = n14022 & n14109;
  assign n14111 = ~n3177 & ~n14110;
  assign n14112 = ~n2980 & n14111;
  assign n14113 = ~n14022 & ~n14109;
  assign n14114 = n13696 & ~n13862;
  assign n14115 = n14114 ^ n13698;
  assign n14116 = n2980 & ~n14115;
  assign n14117 = n14113 & ~n14116;
  assign n14118 = n13702 & ~n13862;
  assign n14119 = n14118 ^ n13704;
  assign n14120 = ~n2782 & ~n14119;
  assign n14121 = n14022 & ~n14120;
  assign n14122 = ~n2980 & n14115;
  assign n14123 = n14121 & ~n14122;
  assign n14124 = n14109 & n14123;
  assign n14125 = ~n3211 & n14115;
  assign n14126 = ~n14120 & ~n14125;
  assign n14127 = ~n14124 & ~n14126;
  assign n14128 = ~n14117 & ~n14127;
  assign n14129 = ~n14112 & n14128;
  assign n14130 = n2782 & n14119;
  assign n14131 = ~n14129 & ~n14130;
  assign n14132 = n14131 ^ n2583;
  assign n14133 = n13708 & ~n13862;
  assign n14134 = n14133 ^ n13710;
  assign n14135 = n14134 ^ n14131;
  assign n14136 = ~n14132 & ~n14135;
  assign n14137 = n14136 ^ n2583;
  assign n14138 = n14137 ^ n2374;
  assign n14139 = n13714 & ~n13862;
  assign n14140 = n14139 ^ n13716;
  assign n14141 = n14140 ^ n14137;
  assign n14142 = n14138 & ~n14141;
  assign n14143 = n14142 ^ n2374;
  assign n14144 = n14143 ^ n2194;
  assign n14145 = n13720 & ~n13862;
  assign n14146 = n14145 ^ n13722;
  assign n14147 = n14146 ^ n14143;
  assign n14148 = ~n14144 & n14147;
  assign n14149 = n14148 ^ n2194;
  assign n14150 = n14149 ^ n2011;
  assign n14151 = n13725 ^ n2194;
  assign n14152 = ~n13862 & ~n14151;
  assign n14153 = n14152 ^ n13571;
  assign n14154 = n14153 ^ n14149;
  assign n14155 = ~n14150 & n14154;
  assign n14156 = n14155 ^ n2011;
  assign n14157 = n14156 ^ n1804;
  assign n14158 = n13725 ^ n13571;
  assign n14159 = ~n14151 & ~n14158;
  assign n14160 = n14159 ^ n2194;
  assign n14161 = n14160 ^ n2011;
  assign n14162 = ~n13862 & ~n14161;
  assign n14163 = n14162 ^ n13728;
  assign n14164 = n14163 ^ n14156;
  assign n14165 = n14157 & n14164;
  assign n14166 = n14165 ^ n1804;
  assign n14167 = n14166 ^ n1621;
  assign n14168 = ~n13742 & ~n13862;
  assign n14169 = n14168 ^ n13745;
  assign n14170 = n14169 ^ n14166;
  assign n14171 = n14167 & ~n14170;
  assign n14172 = n14171 ^ n1621;
  assign n14173 = n14172 ^ n1458;
  assign n14174 = n13749 & ~n13862;
  assign n14175 = n14174 ^ n13752;
  assign n14176 = n14175 ^ n14172;
  assign n14177 = n14173 & n14176;
  assign n14178 = n14177 ^ n1458;
  assign n14179 = n14178 ^ n1299;
  assign n14180 = n13755 ^ n1458;
  assign n14181 = ~n13862 & n14180;
  assign n14182 = n14181 ^ n13567;
  assign n14183 = n14182 ^ n14178;
  assign n14184 = n14179 & ~n14183;
  assign n14185 = n14184 ^ n1299;
  assign n14186 = n14185 ^ n1158;
  assign n14187 = n13758 ^ n1299;
  assign n14188 = ~n13862 & n14187;
  assign n14189 = n14188 ^ n13563;
  assign n14190 = n14189 ^ n14185;
  assign n14191 = n14186 & n14190;
  assign n14192 = n14191 ^ n1158;
  assign n14193 = n14192 ^ n1027;
  assign n14194 = n13762 & ~n13862;
  assign n14195 = n14194 ^ n13764;
  assign n14196 = n14195 ^ n14192;
  assign n14197 = n14193 & ~n14196;
  assign n14198 = n14197 ^ n1027;
  assign n14199 = n14198 ^ n905;
  assign n14200 = n13768 & ~n13862;
  assign n14201 = n14200 ^ n13770;
  assign n14202 = n14201 ^ n14198;
  assign n14203 = n14199 & n14202;
  assign n14204 = n14203 ^ n905;
  assign n14205 = n14204 ^ n803;
  assign n14206 = n13774 & ~n13862;
  assign n14207 = n14206 ^ n13776;
  assign n14208 = n14207 ^ n14204;
  assign n14209 = n14205 & ~n14208;
  assign n14210 = n14209 ^ n803;
  assign n14211 = n14210 ^ n707;
  assign n14212 = n13780 & ~n13862;
  assign n14213 = n14212 ^ n13782;
  assign n14214 = n14213 ^ n14210;
  assign n14215 = ~n14211 & n14214;
  assign n14216 = n14215 ^ n707;
  assign n14217 = n14216 ^ n608;
  assign n14218 = ~n13786 & ~n13862;
  assign n14219 = n14218 ^ n13788;
  assign n14220 = n14219 ^ n14216;
  assign n14221 = ~n14217 & n14220;
  assign n14222 = n14221 ^ n608;
  assign n14223 = n14222 ^ n514;
  assign n14224 = ~n13792 & ~n13862;
  assign n14225 = n14224 ^ n13794;
  assign n14226 = n14225 ^ n14222;
  assign n14227 = n14223 & n14226;
  assign n14228 = n14227 ^ n514;
  assign n14229 = n14228 ^ n436;
  assign n14230 = n13798 & ~n13862;
  assign n14231 = n14230 ^ n13800;
  assign n14232 = n14231 ^ n14228;
  assign n14233 = n14229 & ~n14232;
  assign n14234 = n14233 ^ n436;
  assign n14235 = n14234 ^ n363;
  assign n14236 = n13804 & ~n13862;
  assign n14237 = n14236 ^ n13807;
  assign n14238 = n14237 ^ n14234;
  assign n14239 = n14235 & n14238;
  assign n14240 = n14239 ^ n363;
  assign n14241 = n14240 ^ n300;
  assign n14242 = n13811 & ~n13862;
  assign n14243 = n14242 ^ n13817;
  assign n14244 = n14243 ^ n14240;
  assign n14245 = n14241 & ~n14244;
  assign n14246 = n14245 ^ n300;
  assign n14247 = n14246 ^ n14019;
  assign n14248 = ~n14020 & n14247;
  assign n14249 = n14248 ^ n243;
  assign n14250 = n14249 ^ n14016;
  assign n14251 = n14017 & ~n14250;
  assign n14252 = n14251 ^ n210;
  assign n14253 = n14252 ^ n147;
  assign n14254 = n13833 & ~n13862;
  assign n14255 = n14254 ^ n13836;
  assign n14256 = n14255 ^ n14252;
  assign n14257 = ~n14253 & n14256;
  assign n14258 = n14257 ^ n147;
  assign n14259 = n14258 ^ n132;
  assign n14260 = ~n13840 & ~n13862;
  assign n14261 = n14260 ^ n13846;
  assign n14262 = n14261 ^ n14258;
  assign n14263 = n14259 & n14262;
  assign n14264 = n14263 ^ n132;
  assign n14013 = n13850 & ~n13862;
  assign n14014 = n14013 ^ n13852;
  assign n14265 = n14264 ^ n14014;
  assign n14266 = n14014 ^ n133;
  assign n14267 = n14265 & ~n14266;
  assign n14268 = n14267 ^ n14014;
  assign n14269 = n14012 & n14268;
  assign n14270 = n14008 & ~n14269;
  assign n14271 = n14270 ^ n14028;
  assign n14272 = ~n6181 & n14271;
  assign n14273 = n14002 & ~n14269;
  assign n14274 = n14273 ^ n14004;
  assign n14275 = ~n6479 & ~n14274;
  assign n14276 = ~n14272 & ~n14275;
  assign n14277 = n13915 & ~n14269;
  assign n14278 = n14277 ^ n13917;
  assign n14279 = ~n11820 & n14278;
  assign n14280 = n13870 ^ n13862;
  assign n14281 = ~n14269 & ~n14280;
  assign n14282 = n14281 ^ n13862;
  assign n14283 = n14282 ^ x10;
  assign n14284 = n14283 ^ n13444;
  assign n14285 = ~x6 & ~x7;
  assign n14286 = ~n13862 & n14285;
  assign n14287 = ~x8 & n14286;
  assign n14288 = n13862 & n14285;
  assign n14289 = ~x8 & n14288;
  assign n14290 = n14289 ^ n13862;
  assign n14291 = n14290 ^ n14269;
  assign n14292 = n14291 ^ x9;
  assign n14293 = n14292 ^ n14269;
  assign n14294 = n14293 ^ n14291;
  assign n14295 = ~x8 & ~n14269;
  assign n14296 = n14295 ^ n14291;
  assign n14297 = ~n14294 & ~n14296;
  assign n14298 = n14297 ^ n14292;
  assign n14299 = ~n14287 & ~n14298;
  assign n14300 = n14299 ^ n14283;
  assign n14301 = ~n14284 & n14300;
  assign n14302 = n14301 ^ n13444;
  assign n14303 = n14302 ^ n13031;
  assign n14305 = n13871 ^ n13444;
  assign n14306 = n14305 ^ x10;
  assign n14307 = n14306 ^ n14305;
  assign n14308 = n14305 ^ n13871;
  assign n14309 = n14307 & n14308;
  assign n14310 = n14309 ^ n14305;
  assign n14311 = ~n13862 & ~n14310;
  assign n14312 = n14311 ^ n14305;
  assign n14304 = ~x10 & ~n13862;
  assign n14313 = n14312 ^ n14304;
  assign n14314 = n13870 ^ n13444;
  assign n14315 = n14314 ^ n14312;
  assign n14316 = n14312 ^ n14269;
  assign n14317 = n14312 & ~n14316;
  assign n14318 = n14317 ^ n14312;
  assign n14319 = n14315 & n14318;
  assign n14320 = n14319 ^ n14317;
  assign n14321 = n14320 ^ n14312;
  assign n14322 = n14321 ^ n14269;
  assign n14323 = ~n14313 & ~n14322;
  assign n14324 = n14323 ^ n14304;
  assign n14325 = n14324 ^ x11;
  assign n14326 = n14325 ^ n14302;
  assign n14327 = n14303 & ~n14326;
  assign n14328 = n14327 ^ n13031;
  assign n14329 = n14328 ^ n12617;
  assign n14330 = n13881 & ~n14269;
  assign n14331 = n14330 ^ n13885;
  assign n14332 = n14331 ^ n14328;
  assign n14333 = n14329 & n14332;
  assign n14334 = n14333 ^ n12617;
  assign n14335 = n14334 ^ n12230;
  assign n14336 = n13889 & ~n14269;
  assign n14337 = n14336 ^ n13911;
  assign n14338 = n14337 ^ n14334;
  assign n14339 = n14335 & ~n14338;
  assign n14340 = n14339 ^ n12230;
  assign n14341 = ~n14279 & n14340;
  assign n14342 = n11395 & n11820;
  assign n14343 = n13921 & ~n14269;
  assign n14344 = n14343 ^ n13923;
  assign n14345 = ~n14342 & ~n14344;
  assign n14346 = n14341 & ~n14345;
  assign n14347 = n11395 & ~n14278;
  assign n14348 = n14340 & n14347;
  assign n14349 = n14344 ^ n11395;
  assign n14350 = n11820 & ~n14278;
  assign n14351 = n14350 ^ n14344;
  assign n14352 = n14349 & ~n14351;
  assign n14353 = n14352 ^ n11395;
  assign n14354 = ~n14348 & ~n14353;
  assign n14355 = ~n14346 & n14354;
  assign n14356 = n14355 ^ n10956;
  assign n14357 = n13927 & ~n14269;
  assign n14358 = n14357 ^ n13929;
  assign n14359 = n14358 ^ n14355;
  assign n14360 = ~n14356 & ~n14359;
  assign n14361 = n14360 ^ n10956;
  assign n14362 = n14361 ^ n10585;
  assign n14363 = n13933 & ~n14269;
  assign n14364 = n14363 ^ n13935;
  assign n14365 = n14364 ^ n14361;
  assign n14366 = ~n14362 & ~n14365;
  assign n14367 = n14366 ^ n10585;
  assign n14368 = n14367 ^ n10229;
  assign n14369 = ~n13939 & ~n14269;
  assign n14370 = n14369 ^ n13941;
  assign n14371 = n14370 ^ n14367;
  assign n14372 = ~n14368 & n14371;
  assign n14373 = n14372 ^ n10229;
  assign n14374 = n14373 ^ n9867;
  assign n14375 = ~n13945 & ~n14269;
  assign n14376 = n14375 ^ n13947;
  assign n14377 = n14376 ^ n14373;
  assign n14378 = n14374 & ~n14377;
  assign n14379 = n14378 ^ n9867;
  assign n14380 = n9502 & n14379;
  assign n14381 = n13951 & ~n14269;
  assign n14382 = n14381 ^ n13953;
  assign n14383 = ~n14380 & n14382;
  assign n14384 = n10229 & ~n14367;
  assign n14385 = n14376 & n14384;
  assign n14386 = n14370 ^ n9867;
  assign n14387 = n14370 ^ n10229;
  assign n14388 = n14387 ^ n10229;
  assign n14389 = n14376 ^ n10229;
  assign n14390 = n14388 & ~n14389;
  assign n14391 = n14390 ^ n10229;
  assign n14392 = n14386 & ~n14391;
  assign n14393 = n14392 ^ n9867;
  assign n14394 = ~n14367 & n14393;
  assign n14395 = n14376 ^ n9867;
  assign n14396 = n10229 & n14370;
  assign n14397 = n14396 ^ n9867;
  assign n14398 = n14395 & n14397;
  assign n14399 = n14398 ^ n9867;
  assign n14400 = ~n9502 & ~n14399;
  assign n14401 = ~n14394 & n14400;
  assign n14402 = ~n14385 & n14401;
  assign n14403 = ~n14383 & ~n14402;
  assign n14404 = n14403 ^ n9129;
  assign n14405 = n13957 & ~n14269;
  assign n14406 = n14405 ^ n13959;
  assign n14407 = n14406 ^ n14403;
  assign n14408 = n14404 & ~n14407;
  assign n14409 = n14408 ^ n9129;
  assign n14410 = n14409 ^ n8769;
  assign n14411 = n13963 & ~n14269;
  assign n14412 = n14411 ^ n13965;
  assign n14413 = n14412 ^ n14409;
  assign n14414 = n14410 & n14413;
  assign n14415 = n14414 ^ n8769;
  assign n14416 = n14415 ^ n8422;
  assign n14417 = n13969 & ~n14269;
  assign n14418 = n14417 ^ n13972;
  assign n14419 = n14418 ^ n14415;
  assign n14420 = n14416 & ~n14419;
  assign n14421 = n14420 ^ n8422;
  assign n14422 = n14421 ^ n8083;
  assign n14423 = n13976 & ~n14269;
  assign n14424 = n14423 ^ n13979;
  assign n14425 = n14424 ^ n14421;
  assign n14426 = n14422 & n14425;
  assign n14427 = n14426 ^ n8083;
  assign n14428 = n14427 ^ n7777;
  assign n14429 = n13982 ^ n8083;
  assign n14430 = ~n14269 & n14429;
  assign n14431 = n14430 ^ n13867;
  assign n14432 = n14431 ^ n14427;
  assign n14433 = n14428 & ~n14432;
  assign n14434 = n14433 ^ n7777;
  assign n14435 = n14434 ^ n7463;
  assign n14436 = n13982 ^ n13867;
  assign n14437 = n14429 & ~n14436;
  assign n14438 = n14437 ^ n8083;
  assign n14439 = n14438 ^ n7777;
  assign n14440 = ~n14269 & n14439;
  assign n14441 = n14440 ^ n13864;
  assign n14442 = n14441 ^ n14434;
  assign n14443 = n14435 & ~n14442;
  assign n14444 = n14443 ^ n7463;
  assign n14445 = n14444 ^ n7135;
  assign n14446 = ~n13990 & ~n14269;
  assign n14447 = n14446 ^ n13992;
  assign n14448 = n14447 ^ n14444;
  assign n14449 = n14445 & ~n14448;
  assign n14450 = n14449 ^ n7135;
  assign n14451 = n14450 ^ n6802;
  assign n14452 = n13996 & ~n14269;
  assign n14453 = n14452 ^ n13998;
  assign n14454 = n14453 ^ n14450;
  assign n14455 = n14451 & n14454;
  assign n14456 = n14455 ^ n6802;
  assign n14457 = n14276 & n14456;
  assign n14458 = n14271 ^ n6181;
  assign n14459 = n6479 & n14274;
  assign n14460 = n14459 ^ n14271;
  assign n14461 = ~n14458 & n14460;
  assign n14462 = n14461 ^ n6181;
  assign n14463 = ~n14457 & ~n14462;
  assign n14464 = n14463 ^ n5905;
  assign n14465 = n14259 & ~n14269;
  assign n14466 = n14465 ^ n14261;
  assign n14467 = ~n133 & ~n14466;
  assign n14468 = n14241 & ~n14269;
  assign n14469 = n14468 ^ n14243;
  assign n14470 = ~n243 & ~n14469;
  assign n14471 = n14173 & ~n14269;
  assign n14472 = n14471 ^ n14175;
  assign n14473 = n14472 ^ n1299;
  assign n14474 = n14167 & ~n14269;
  assign n14475 = n14474 ^ n14169;
  assign n14476 = n14475 ^ n1458;
  assign n14477 = n14032 & ~n14269;
  assign n14478 = n14477 ^ n14034;
  assign n14479 = n14478 ^ n14463;
  assign n14480 = ~n14464 & n14479;
  assign n14481 = n14480 ^ n5905;
  assign n14482 = n14481 ^ n5625;
  assign n14483 = n14038 & ~n14269;
  assign n14484 = n14483 ^ n14040;
  assign n14485 = n14484 ^ n14481;
  assign n14486 = n14482 & n14485;
  assign n14487 = n14486 ^ n5625;
  assign n14488 = n14487 ^ n5363;
  assign n14489 = n14044 & ~n14269;
  assign n14490 = n14489 ^ n14046;
  assign n14491 = n14490 ^ n14487;
  assign n14492 = n14488 & ~n14491;
  assign n14493 = n14492 ^ n5363;
  assign n14494 = n14493 ^ n5108;
  assign n14495 = n14049 ^ n5363;
  assign n14496 = ~n14269 & n14495;
  assign n14497 = n14496 ^ n14025;
  assign n14498 = n14497 ^ n14493;
  assign n14499 = n14494 & n14498;
  assign n14500 = n14499 ^ n5108;
  assign n14501 = n14500 ^ n4851;
  assign n14502 = ~n14050 & ~n14060;
  assign n14503 = n14502 ^ n5108;
  assign n14504 = ~n14269 & ~n14503;
  assign n14505 = n14504 ^ n14054;
  assign n14506 = n14505 ^ n14500;
  assign n14507 = n14501 & ~n14506;
  assign n14508 = n14507 ^ n4851;
  assign n14509 = n14508 ^ n4606;
  assign n14510 = ~n14066 & ~n14269;
  assign n14511 = n14510 ^ n14068;
  assign n14512 = n14511 ^ n14508;
  assign n14513 = n14509 & n14512;
  assign n14514 = n14513 ^ n4606;
  assign n14515 = n14514 ^ n4362;
  assign n14516 = n14072 & ~n14269;
  assign n14517 = n14516 ^ n14074;
  assign n14518 = n14517 ^ n14514;
  assign n14519 = n14515 & ~n14518;
  assign n14520 = n14519 ^ n4362;
  assign n14521 = n14520 ^ n4133;
  assign n14522 = n14078 & ~n14269;
  assign n14523 = n14522 ^ n14080;
  assign n14524 = n14523 ^ n14520;
  assign n14525 = n14521 & n14524;
  assign n14526 = n14525 ^ n4133;
  assign n14527 = n14526 ^ n3882;
  assign n14528 = n14084 & ~n14269;
  assign n14529 = n14528 ^ n14086;
  assign n14530 = n14529 ^ n14526;
  assign n14531 = n14527 & ~n14530;
  assign n14532 = n14531 ^ n3882;
  assign n14533 = n14532 ^ n3634;
  assign n14534 = n14090 & ~n14269;
  assign n14535 = n14534 ^ n14093;
  assign n14536 = n14535 ^ n14532;
  assign n14537 = ~n14533 & n14536;
  assign n14538 = n14537 ^ n3634;
  assign n14539 = n14538 ^ n3397;
  assign n14540 = ~n14097 & ~n14269;
  assign n14541 = n14540 ^ n14100;
  assign n14542 = n14541 ^ n14538;
  assign n14543 = ~n14539 & n14542;
  assign n14544 = n14543 ^ n3397;
  assign n14545 = n14544 ^ n3177;
  assign n14546 = ~n14104 & ~n14269;
  assign n14547 = n14546 ^ n14106;
  assign n14548 = n14547 ^ n14544;
  assign n14549 = n14545 & ~n14548;
  assign n14550 = n14549 ^ n3177;
  assign n14551 = n14550 ^ n2980;
  assign n14552 = n14109 ^ n3177;
  assign n14553 = ~n14269 & n14552;
  assign n14554 = n14553 ^ n14022;
  assign n14555 = n14554 ^ n14550;
  assign n14556 = n14551 & ~n14555;
  assign n14557 = n14556 ^ n2980;
  assign n14558 = n14557 ^ n2782;
  assign n14559 = ~n14111 & ~n14113;
  assign n14560 = n14559 ^ n2980;
  assign n14561 = ~n14269 & n14560;
  assign n14562 = n14561 ^ n14115;
  assign n14563 = n14562 ^ n14557;
  assign n14564 = n14558 & n14563;
  assign n14565 = n14564 ^ n2782;
  assign n14566 = n14565 ^ n2583;
  assign n14567 = n14115 ^ n2980;
  assign n14568 = n14559 ^ n14115;
  assign n14569 = ~n14567 & n14568;
  assign n14570 = n14569 ^ n2980;
  assign n14571 = n14570 ^ n2782;
  assign n14572 = ~n14269 & n14571;
  assign n14573 = n14572 ^ n14119;
  assign n14574 = n14573 ^ n14565;
  assign n14575 = n14566 & ~n14574;
  assign n14576 = n14575 ^ n2583;
  assign n14577 = n14576 ^ n2374;
  assign n14578 = ~n14132 & ~n14269;
  assign n14579 = n14578 ^ n14134;
  assign n14580 = n14579 ^ n14576;
  assign n14581 = n14577 & n14580;
  assign n14582 = n14581 ^ n2374;
  assign n14583 = n14582 ^ n2194;
  assign n14584 = n14138 & ~n14269;
  assign n14585 = n14584 ^ n14140;
  assign n14586 = n14585 ^ n14582;
  assign n14587 = ~n14583 & ~n14586;
  assign n14588 = n14587 ^ n2194;
  assign n14589 = n14588 ^ n2011;
  assign n14590 = ~n14144 & ~n14269;
  assign n14591 = n14590 ^ n14146;
  assign n14592 = n14591 ^ n14588;
  assign n14593 = ~n14589 & ~n14592;
  assign n14594 = n14593 ^ n2011;
  assign n14595 = n14594 ^ n1804;
  assign n14596 = ~n14150 & ~n14269;
  assign n14597 = n14596 ^ n14153;
  assign n14598 = n14597 ^ n14594;
  assign n14599 = n14595 & ~n14598;
  assign n14600 = n14599 ^ n1804;
  assign n14601 = n14600 ^ n1621;
  assign n14602 = n14157 & ~n14269;
  assign n14603 = n14602 ^ n14163;
  assign n14604 = n14603 ^ n14600;
  assign n14605 = n14601 & n14604;
  assign n14606 = n14605 ^ n1621;
  assign n14607 = n14606 ^ n14475;
  assign n14608 = n14476 & ~n14607;
  assign n14609 = n14608 ^ n1458;
  assign n14610 = n14609 ^ n14472;
  assign n14611 = ~n14473 & n14610;
  assign n14612 = n14611 ^ n1299;
  assign n14613 = n14612 ^ n1158;
  assign n14614 = n14179 & ~n14269;
  assign n14615 = n14614 ^ n14182;
  assign n14616 = n14615 ^ n14612;
  assign n14617 = n14613 & ~n14616;
  assign n14618 = n14617 ^ n1158;
  assign n14619 = n14618 ^ n1027;
  assign n14620 = n14186 & ~n14269;
  assign n14621 = n14620 ^ n14189;
  assign n14622 = n14621 ^ n14618;
  assign n14623 = n14619 & n14622;
  assign n14624 = n14623 ^ n1027;
  assign n14625 = n14624 ^ n905;
  assign n14626 = n14193 & ~n14269;
  assign n14627 = n14626 ^ n14195;
  assign n14628 = n14627 ^ n14624;
  assign n14629 = n14625 & ~n14628;
  assign n14630 = n14629 ^ n905;
  assign n14631 = n14630 ^ n803;
  assign n14632 = n14199 & ~n14269;
  assign n14633 = n14632 ^ n14201;
  assign n14634 = n14633 ^ n14630;
  assign n14635 = n14631 & n14634;
  assign n14636 = n14635 ^ n803;
  assign n14637 = n14636 ^ n707;
  assign n14638 = n14205 & ~n14269;
  assign n14639 = n14638 ^ n14207;
  assign n14640 = n14639 ^ n14636;
  assign n14641 = ~n14637 & ~n14640;
  assign n14642 = n14641 ^ n707;
  assign n14643 = n14642 ^ n608;
  assign n14644 = ~n14211 & ~n14269;
  assign n14645 = n14644 ^ n14213;
  assign n14646 = n14645 ^ n14642;
  assign n14647 = ~n14643 & ~n14646;
  assign n14648 = n14647 ^ n608;
  assign n14649 = n14648 ^ n514;
  assign n14650 = ~n14217 & ~n14269;
  assign n14651 = n14650 ^ n14219;
  assign n14652 = n14651 ^ n14648;
  assign n14653 = n14649 & ~n14652;
  assign n14654 = n14653 ^ n514;
  assign n14655 = n14654 ^ n436;
  assign n14656 = n14223 & ~n14269;
  assign n14657 = n14656 ^ n14225;
  assign n14658 = n14657 ^ n14654;
  assign n14659 = n14655 & n14658;
  assign n14660 = n14659 ^ n436;
  assign n14661 = n14660 ^ n363;
  assign n14662 = n14229 & ~n14269;
  assign n14663 = n14662 ^ n14231;
  assign n14664 = n14663 ^ n14660;
  assign n14665 = n14661 & ~n14664;
  assign n14666 = n14665 ^ n363;
  assign n14667 = n14666 ^ n300;
  assign n14668 = n14235 & ~n14269;
  assign n14669 = n14668 ^ n14237;
  assign n14670 = n14669 ^ n14666;
  assign n14671 = n14667 & n14670;
  assign n14672 = n14671 ^ n300;
  assign n14673 = ~n14470 & n14672;
  assign n14674 = n210 & n243;
  assign n14675 = n14246 ^ n243;
  assign n14676 = ~n14269 & n14675;
  assign n14677 = n14676 ^ n14019;
  assign n14678 = ~n14674 & n14677;
  assign n14679 = n14673 & ~n14678;
  assign n14680 = n210 & n14469;
  assign n14681 = n14672 & n14680;
  assign n14682 = n14677 ^ n210;
  assign n14683 = n243 & n14469;
  assign n14684 = n14683 ^ n14677;
  assign n14685 = ~n14682 & n14684;
  assign n14686 = n14685 ^ n210;
  assign n14687 = ~n14681 & ~n14686;
  assign n14688 = ~n14679 & n14687;
  assign n14689 = n14688 ^ n147;
  assign n14690 = n14249 ^ n210;
  assign n14691 = ~n14269 & n14690;
  assign n14692 = n14691 ^ n14016;
  assign n14693 = n14692 ^ n14688;
  assign n14694 = n14689 & n14693;
  assign n14695 = n14694 ^ n147;
  assign n14696 = n14695 ^ n132;
  assign n14697 = ~n14253 & ~n14269;
  assign n14698 = n14697 ^ n14255;
  assign n14699 = n14698 ^ n14695;
  assign n14700 = n14696 & ~n14699;
  assign n14701 = n14700 ^ n132;
  assign n14702 = ~n14467 & ~n14701;
  assign n14703 = ~n14012 & n14014;
  assign n14704 = n14703 ^ n14014;
  assign n14708 = n14265 ^ n14014;
  assign n14709 = ~n14704 & ~n14708;
  assign n14710 = n14709 ^ n14014;
  assign n14705 = n14264 & ~n14704;
  assign n14706 = n14705 ^ n14014;
  assign n14707 = ~n14466 & n14706;
  assign n14711 = n14710 ^ n14707;
  assign n14712 = ~n133 & n14711;
  assign n14713 = n14712 ^ n14707;
  assign n14714 = ~n14702 & n14713;
  assign n14715 = ~n14464 & ~n14714;
  assign n14716 = n14715 ^ n14478;
  assign n14717 = n14716 ^ n5625;
  assign n14718 = n14456 ^ n6479;
  assign n14719 = n14456 ^ n14274;
  assign n14720 = n14718 & ~n14719;
  assign n14721 = n14720 ^ n6479;
  assign n14722 = n14721 ^ n6181;
  assign n14723 = ~n14714 & n14722;
  assign n14724 = n14723 ^ n14271;
  assign n14725 = n14724 ^ n5905;
  assign n14726 = ~n14356 & ~n14714;
  assign n14727 = n14726 ^ n14358;
  assign n14728 = ~n14341 & ~n14350;
  assign n14729 = n14728 ^ n11395;
  assign n14730 = ~n14714 & ~n14729;
  assign n14731 = n14730 ^ n14344;
  assign n14732 = n14731 ^ n10956;
  assign n14733 = n14340 ^ n11820;
  assign n14734 = ~n14714 & n14733;
  assign n14735 = n14734 ^ n14278;
  assign n14736 = n14735 ^ n11395;
  assign n14737 = ~x4 & ~x5;
  assign n14738 = ~x6 & n14737;
  assign n14739 = n14269 & ~n14738;
  assign n14740 = n14714 ^ x7;
  assign n14741 = ~n14739 & n14740;
  assign n14743 = ~n14269 & n14737;
  assign n14742 = ~x7 & ~n14714;
  assign n14744 = n14743 ^ n14742;
  assign n14745 = ~x6 & n14744;
  assign n14746 = n14745 ^ n14742;
  assign n14747 = ~n14741 & ~n14746;
  assign n14748 = n14747 ^ n13862;
  assign n14749 = n14285 ^ n14269;
  assign n14750 = ~n14714 & ~n14749;
  assign n14751 = n14750 ^ n14269;
  assign n14752 = n14751 ^ x8;
  assign n14753 = n14752 ^ n14747;
  assign n14754 = n14748 & n14753;
  assign n14755 = n14754 ^ n13862;
  assign n14756 = n14755 ^ n13444;
  assign n14757 = n14269 ^ n13862;
  assign n14758 = n14757 ^ n14269;
  assign n14759 = n14758 ^ n14757;
  assign n14760 = n14757 ^ n14285;
  assign n14761 = n14759 & n14760;
  assign n14762 = n14761 ^ n14757;
  assign n14763 = ~x8 & n14762;
  assign n14764 = n14763 ^ n14757;
  assign n14765 = n14764 ^ n14295;
  assign n14766 = n14285 ^ n13862;
  assign n14767 = n14766 ^ n14764;
  assign n14768 = n14764 ^ n14714;
  assign n14769 = ~n14764 & n14768;
  assign n14770 = n14769 ^ n14764;
  assign n14771 = ~n14767 & ~n14770;
  assign n14772 = n14771 ^ n14769;
  assign n14773 = n14772 ^ n14764;
  assign n14774 = n14773 ^ n14714;
  assign n14775 = n14765 & n14774;
  assign n14776 = n14775 ^ n14295;
  assign n14777 = n14776 ^ x9;
  assign n14778 = n14777 ^ n14755;
  assign n14779 = n14756 & ~n14778;
  assign n14780 = n14779 ^ n13444;
  assign n14781 = n14780 ^ n13031;
  assign n14782 = n14299 ^ n13444;
  assign n14783 = ~n14714 & n14782;
  assign n14784 = n14783 ^ n14283;
  assign n14785 = n14784 ^ n14780;
  assign n14786 = n14781 & n14785;
  assign n14787 = n14786 ^ n13031;
  assign n14788 = n14787 ^ n12617;
  assign n14789 = n14303 & ~n14714;
  assign n14790 = n14789 ^ n14325;
  assign n14791 = n14790 ^ n14787;
  assign n14792 = n14788 & ~n14791;
  assign n14793 = n14792 ^ n12617;
  assign n14794 = n14793 ^ n12230;
  assign n14795 = n14329 & ~n14714;
  assign n14796 = n14795 ^ n14331;
  assign n14797 = n14796 ^ n14793;
  assign n14798 = n14794 & n14797;
  assign n14799 = n14798 ^ n12230;
  assign n14800 = n14799 ^ n11820;
  assign n14801 = n14335 & ~n14714;
  assign n14802 = n14801 ^ n14337;
  assign n14803 = n14802 ^ n14799;
  assign n14804 = n14800 & ~n14803;
  assign n14805 = n14804 ^ n11820;
  assign n14806 = n14805 ^ n14735;
  assign n14807 = ~n14736 & n14806;
  assign n14808 = n14807 ^ n11395;
  assign n14809 = n14808 ^ n14731;
  assign n14810 = n14732 & ~n14809;
  assign n14811 = n14810 ^ n10956;
  assign n14812 = ~n14727 & n14811;
  assign n14813 = ~n10585 & n14811;
  assign n14814 = ~n14812 & ~n14813;
  assign n14815 = n10229 & ~n10585;
  assign n14816 = ~n14362 & ~n14714;
  assign n14817 = n14816 ^ n14364;
  assign n14818 = ~n14815 & ~n14817;
  assign n14819 = ~n14814 & ~n14818;
  assign n14820 = ~n14727 & n14815;
  assign n14821 = ~n14817 & ~n14820;
  assign n14822 = ~n14812 & n14821;
  assign n14823 = ~n10585 & ~n14727;
  assign n14824 = n14817 & n14823;
  assign n14825 = ~n10229 & ~n14824;
  assign n14826 = ~n14822 & ~n14825;
  assign n14827 = ~n14819 & ~n14826;
  assign n14828 = n14827 ^ n9867;
  assign n14829 = ~n14368 & ~n14714;
  assign n14830 = n14829 ^ n14370;
  assign n14831 = n14830 ^ n14827;
  assign n14832 = ~n14828 & n14831;
  assign n14833 = n14832 ^ n9867;
  assign n14834 = n14833 ^ n9502;
  assign n14835 = n14374 & ~n14714;
  assign n14836 = n14835 ^ n14376;
  assign n14837 = n14836 ^ n14833;
  assign n14838 = n14834 & ~n14837;
  assign n14839 = n14838 ^ n9502;
  assign n14840 = n14839 ^ n9129;
  assign n14841 = n14379 ^ n9502;
  assign n14842 = ~n14714 & n14841;
  assign n14843 = n14842 ^ n14382;
  assign n14844 = n14843 ^ n14839;
  assign n14845 = n14840 & n14844;
  assign n14846 = n14845 ^ n9129;
  assign n14847 = n14846 ^ n8769;
  assign n14848 = n14404 & ~n14714;
  assign n14849 = n14848 ^ n14406;
  assign n14850 = n14849 ^ n14846;
  assign n14851 = n14847 & ~n14850;
  assign n14852 = n14851 ^ n8769;
  assign n14853 = n14852 ^ n8422;
  assign n14854 = n14410 & ~n14714;
  assign n14855 = n14854 ^ n14412;
  assign n14856 = n14855 ^ n14852;
  assign n14857 = n14853 & n14856;
  assign n14858 = n14857 ^ n8422;
  assign n14859 = n14858 ^ n8083;
  assign n14860 = n14416 & ~n14714;
  assign n14861 = n14860 ^ n14418;
  assign n14862 = n14861 ^ n14858;
  assign n14863 = n14859 & ~n14862;
  assign n14864 = n14863 ^ n8083;
  assign n14865 = n14864 ^ n7777;
  assign n14866 = n14422 & ~n14714;
  assign n14867 = n14866 ^ n14424;
  assign n14868 = n14867 ^ n14864;
  assign n14869 = n14865 & n14868;
  assign n14870 = n14869 ^ n7777;
  assign n14871 = n14870 ^ n7463;
  assign n14872 = n14428 & ~n14714;
  assign n14873 = n14872 ^ n14431;
  assign n14874 = n14873 ^ n14870;
  assign n14875 = n14871 & ~n14874;
  assign n14876 = n14875 ^ n7463;
  assign n14877 = n14876 ^ n7135;
  assign n14878 = n14435 & ~n14714;
  assign n14879 = n14878 ^ n14441;
  assign n14880 = n14879 ^ n14876;
  assign n14881 = n14877 & ~n14880;
  assign n14882 = n14881 ^ n7135;
  assign n14883 = n14882 ^ n6802;
  assign n14884 = n14445 & ~n14714;
  assign n14885 = n14884 ^ n14447;
  assign n14886 = n14885 ^ n14882;
  assign n14887 = n14883 & ~n14886;
  assign n14888 = n14887 ^ n6802;
  assign n14889 = n14888 ^ n6479;
  assign n14890 = n14451 & ~n14714;
  assign n14891 = n14890 ^ n14453;
  assign n14892 = n14891 ^ n14888;
  assign n14893 = n14889 & n14892;
  assign n14894 = n14893 ^ n6479;
  assign n14895 = n14894 ^ n6181;
  assign n14896 = ~n14714 & n14718;
  assign n14897 = n14896 ^ n14274;
  assign n14898 = n14897 ^ n14894;
  assign n14899 = n14895 & ~n14898;
  assign n14900 = n14899 ^ n6181;
  assign n14901 = n14900 ^ n14724;
  assign n14902 = ~n14725 & n14901;
  assign n14903 = n14902 ^ n5905;
  assign n14904 = n14903 ^ n14716;
  assign n14905 = n14717 & ~n14904;
  assign n14906 = n14905 ^ n5625;
  assign n14907 = n14906 ^ n5363;
  assign n14908 = n14482 & ~n14714;
  assign n14909 = n14908 ^ n14484;
  assign n14910 = n14909 ^ n14906;
  assign n14911 = n14907 & n14910;
  assign n14912 = n14911 ^ n5363;
  assign n14913 = n14912 ^ n5108;
  assign n14914 = n14488 & ~n14714;
  assign n14915 = n14914 ^ n14490;
  assign n14916 = n14915 ^ n14912;
  assign n14917 = n14913 & ~n14916;
  assign n14918 = n14917 ^ n5108;
  assign n14919 = n14918 ^ n4851;
  assign n14920 = n14494 & ~n14714;
  assign n14921 = n14920 ^ n14497;
  assign n14922 = n14921 ^ n14918;
  assign n14923 = n14919 & n14922;
  assign n14924 = n14923 ^ n4851;
  assign n14925 = n14924 ^ n4606;
  assign n14926 = n14501 & ~n14714;
  assign n14927 = n14926 ^ n14505;
  assign n14928 = n14927 ^ n14924;
  assign n14929 = n14925 & ~n14928;
  assign n14930 = n14929 ^ n4606;
  assign n14931 = n14930 ^ n4362;
  assign n14932 = n14509 & ~n14714;
  assign n14933 = n14932 ^ n14511;
  assign n14934 = n14933 ^ n14930;
  assign n14935 = n14931 & n14934;
  assign n14936 = n14935 ^ n4362;
  assign n14937 = n14936 ^ n4133;
  assign n14938 = n14515 & ~n14714;
  assign n14939 = n14938 ^ n14517;
  assign n14940 = n14939 ^ n14936;
  assign n14941 = n14937 & ~n14940;
  assign n14942 = n14941 ^ n4133;
  assign n14943 = n14942 ^ n3882;
  assign n14944 = n14521 & ~n14714;
  assign n14945 = n14944 ^ n14523;
  assign n14946 = n14945 ^ n14942;
  assign n14947 = n14943 & n14946;
  assign n14948 = n14947 ^ n3882;
  assign n14949 = n14948 ^ n3634;
  assign n14950 = n14527 & ~n14714;
  assign n14951 = n14950 ^ n14529;
  assign n14952 = n14951 ^ n14948;
  assign n14953 = ~n14949 & ~n14952;
  assign n14954 = n14953 ^ n3634;
  assign n14955 = n14954 ^ n3397;
  assign n14956 = ~n14533 & ~n14714;
  assign n14957 = n14956 ^ n14535;
  assign n14958 = n14957 ^ n14954;
  assign n14959 = ~n14955 & ~n14958;
  assign n14960 = n14959 ^ n3397;
  assign n14961 = n14960 ^ n3177;
  assign n14962 = ~n14539 & ~n14714;
  assign n14963 = n14962 ^ n14541;
  assign n14964 = n14963 ^ n14960;
  assign n14965 = n14961 & ~n14964;
  assign n14966 = n14965 ^ n3177;
  assign n14967 = n14966 ^ n2980;
  assign n14968 = n14545 & ~n14714;
  assign n14969 = n14968 ^ n14547;
  assign n14970 = n14969 ^ n14966;
  assign n14971 = n14967 & ~n14970;
  assign n14972 = n14971 ^ n2980;
  assign n14973 = n14972 ^ n2782;
  assign n14974 = n14551 & ~n14714;
  assign n14975 = n14974 ^ n14554;
  assign n14976 = n14975 ^ n14972;
  assign n14977 = n14973 & ~n14976;
  assign n14978 = n14977 ^ n2782;
  assign n14979 = n14978 ^ n2583;
  assign n14980 = n14558 & ~n14714;
  assign n14981 = n14980 ^ n14562;
  assign n14982 = n14981 ^ n14978;
  assign n14983 = n14979 & n14982;
  assign n14984 = n14983 ^ n2583;
  assign n14985 = n14984 ^ n2374;
  assign n14986 = n14566 & ~n14714;
  assign n14987 = n14986 ^ n14573;
  assign n14988 = n14987 ^ n14984;
  assign n14989 = n14985 & ~n14988;
  assign n14990 = n14989 ^ n2374;
  assign n14991 = n14990 ^ n2194;
  assign n14992 = n14577 & ~n14714;
  assign n14993 = n14992 ^ n14579;
  assign n14994 = n14993 ^ n14990;
  assign n14995 = ~n14991 & n14994;
  assign n14996 = n14995 ^ n2194;
  assign n14997 = n14996 ^ n2011;
  assign n14998 = ~n14583 & ~n14714;
  assign n14999 = n14998 ^ n14585;
  assign n15000 = n14999 ^ n14996;
  assign n15001 = ~n14997 & n15000;
  assign n15002 = n15001 ^ n2011;
  assign n15003 = n15002 ^ n1804;
  assign n15004 = ~n14589 & ~n14714;
  assign n15005 = n15004 ^ n14591;
  assign n15006 = n15005 ^ n15002;
  assign n15007 = n15003 & n15006;
  assign n15008 = n15007 ^ n1804;
  assign n15009 = n15008 ^ n1621;
  assign n15010 = n14595 & ~n14714;
  assign n15011 = n15010 ^ n14597;
  assign n15012 = n15011 ^ n15008;
  assign n15013 = n15009 & ~n15012;
  assign n15014 = n15013 ^ n1621;
  assign n15015 = n15014 ^ n1458;
  assign n15016 = n14601 & ~n14714;
  assign n15017 = n15016 ^ n14603;
  assign n15018 = n15017 ^ n15014;
  assign n15019 = n15015 & n15018;
  assign n15020 = n15019 ^ n1458;
  assign n15021 = n15020 ^ n1299;
  assign n15022 = n14606 ^ n1458;
  assign n15023 = ~n14714 & n15022;
  assign n15024 = n15023 ^ n14475;
  assign n15025 = n15024 ^ n15020;
  assign n15026 = n15021 & ~n15025;
  assign n15027 = n15026 ^ n1299;
  assign n15028 = n15027 ^ n1158;
  assign n15029 = n14609 ^ n1299;
  assign n15030 = ~n14714 & n15029;
  assign n15031 = n15030 ^ n14472;
  assign n15032 = n15031 ^ n15027;
  assign n15033 = n15028 & n15032;
  assign n15034 = n15033 ^ n1158;
  assign n15035 = n15034 ^ n1027;
  assign n15036 = n14613 & ~n14714;
  assign n15037 = n15036 ^ n14615;
  assign n15038 = n15037 ^ n15034;
  assign n15039 = n15035 & ~n15038;
  assign n15040 = n15039 ^ n1027;
  assign n15041 = n15040 ^ n905;
  assign n15042 = n14619 & ~n14714;
  assign n15043 = n15042 ^ n14621;
  assign n15044 = n15043 ^ n15040;
  assign n15045 = n15041 & n15044;
  assign n15046 = n15045 ^ n905;
  assign n15047 = n15046 ^ n803;
  assign n15048 = n14625 & ~n14714;
  assign n15049 = n15048 ^ n14627;
  assign n15050 = n15049 ^ n15046;
  assign n15051 = n15047 & ~n15050;
  assign n15052 = n15051 ^ n803;
  assign n15053 = n15052 ^ n707;
  assign n15054 = n14631 & ~n14714;
  assign n15055 = n15054 ^ n14633;
  assign n15056 = n15055 ^ n15052;
  assign n15057 = ~n15053 & n15056;
  assign n15058 = n15057 ^ n707;
  assign n15059 = n15058 ^ n608;
  assign n15060 = ~n14637 & ~n14714;
  assign n15061 = n15060 ^ n14639;
  assign n15062 = n15061 ^ n15058;
  assign n15063 = ~n15059 & n15062;
  assign n15064 = n15063 ^ n608;
  assign n15065 = n15064 ^ n514;
  assign n15066 = ~n14643 & ~n14714;
  assign n15067 = n15066 ^ n14645;
  assign n15068 = n15067 ^ n15064;
  assign n15069 = n15065 & n15068;
  assign n15070 = n15069 ^ n514;
  assign n15071 = n15070 ^ n436;
  assign n15072 = n14649 & ~n14714;
  assign n15073 = n15072 ^ n14651;
  assign n15074 = n15073 ^ n15070;
  assign n15075 = n15071 & ~n15074;
  assign n15076 = n15075 ^ n436;
  assign n15077 = n15076 ^ n363;
  assign n15078 = n14655 & ~n14714;
  assign n15079 = n15078 ^ n14657;
  assign n15080 = n15079 ^ n15076;
  assign n15081 = n15077 & n15080;
  assign n15082 = n15081 ^ n363;
  assign n15083 = n15082 ^ n300;
  assign n15084 = n14661 & ~n14714;
  assign n15085 = n15084 ^ n14663;
  assign n15086 = n15085 ^ n15082;
  assign n15087 = n15083 & ~n15086;
  assign n15088 = n15087 ^ n300;
  assign n15089 = n15088 ^ n243;
  assign n15090 = n14667 & ~n14714;
  assign n15091 = n15090 ^ n14669;
  assign n15092 = n15091 ^ n15088;
  assign n15093 = n15089 & n15092;
  assign n15094 = n15093 ^ n243;
  assign n15095 = n15094 ^ n210;
  assign n15096 = n14696 & ~n14714;
  assign n15097 = n15096 ^ n14698;
  assign n15098 = n14466 & ~n14701;
  assign n15099 = n15097 & ~n15098;
  assign n15100 = n133 & ~n15099;
  assign n15108 = ~n133 & n14701;
  assign n15101 = n14701 ^ n133;
  assign n15102 = n14710 ^ n14706;
  assign n15103 = n14710 ^ n14701;
  assign n15104 = n15103 ^ n14710;
  assign n15105 = n15102 & n15104;
  assign n15106 = n15105 ^ n14710;
  assign n15107 = ~n15101 & ~n15106;
  assign n15109 = n15108 ^ n15107;
  assign n15110 = ~n14466 & n15109;
  assign n15111 = n15110 ^ n15108;
  assign n15112 = ~n15100 & ~n15111;
  assign n15113 = n14672 ^ n243;
  assign n15114 = ~n14714 & n15113;
  assign n15115 = n15114 ^ n14469;
  assign n15116 = n15115 ^ n15094;
  assign n15117 = n15095 & ~n15116;
  assign n15118 = n15117 ^ n210;
  assign n15119 = n15118 ^ n147;
  assign n15120 = ~n14673 & ~n14683;
  assign n15121 = n15120 ^ n210;
  assign n15122 = ~n14714 & ~n15121;
  assign n15123 = n15122 ^ n14677;
  assign n15124 = n15123 ^ n15118;
  assign n15125 = ~n15119 & n15124;
  assign n15126 = n15125 ^ n147;
  assign n15127 = n15126 ^ n132;
  assign n15128 = n14689 & ~n14714;
  assign n15129 = n15128 ^ n14692;
  assign n15130 = n15129 ^ n15126;
  assign n15131 = n15127 & n15130;
  assign n15132 = n15131 ^ n132;
  assign n15133 = n15097 & ~n15132;
  assign n15134 = ~n133 & n15133;
  assign n15135 = n15134 ^ n15132;
  assign n15136 = n15112 & n15135;
  assign n15137 = n15095 & ~n15136;
  assign n15138 = n15137 ^ n15115;
  assign n15139 = n15138 ^ n147;
  assign n15140 = n15089 & ~n15136;
  assign n15141 = n15140 ^ n15091;
  assign n15142 = n15141 ^ n210;
  assign n15143 = n14925 & ~n15136;
  assign n15144 = n15143 ^ n14927;
  assign n15145 = ~n4362 & ~n15144;
  assign n15146 = n14931 & ~n15136;
  assign n15147 = n15146 ^ n14933;
  assign n15148 = ~n4133 & n15147;
  assign n15149 = ~n15145 & ~n15148;
  assign n15150 = n14756 & ~n15136;
  assign n15151 = n15150 ^ n14777;
  assign n15152 = n15151 ^ n13031;
  assign n15153 = n14748 & ~n15136;
  assign n15154 = n15153 ^ n14752;
  assign n15155 = n15154 ^ n13444;
  assign n15156 = n14737 ^ n14714;
  assign n15157 = ~n15136 & ~n15156;
  assign n15158 = n15157 ^ n14714;
  assign n15159 = n15158 ^ x6;
  assign n15160 = n15159 ^ n14269;
  assign n15161 = ~x2 & ~x3;
  assign n15162 = ~n14714 & n15161;
  assign n15163 = ~x4 & n15162;
  assign n15164 = ~n14737 & ~n15136;
  assign n15165 = n15164 ^ x5;
  assign n15166 = n15164 ^ n15136;
  assign n15167 = n14714 & ~n15161;
  assign n15168 = x4 & n14714;
  assign n15169 = ~n15167 & ~n15168;
  assign n15170 = n15169 ^ n15136;
  assign n15171 = n15170 ^ n15136;
  assign n15172 = n15166 & ~n15171;
  assign n15173 = n15172 ^ n15136;
  assign n15174 = ~n15165 & ~n15173;
  assign n15175 = n15174 ^ x5;
  assign n15176 = ~n15163 & n15175;
  assign n15177 = n15176 ^ n15159;
  assign n15178 = ~n15160 & n15177;
  assign n15179 = n15178 ^ n14269;
  assign n15180 = n15179 ^ n13862;
  assign n15182 = n14738 ^ n14269;
  assign n15183 = n15182 ^ x6;
  assign n15184 = n15183 ^ n15182;
  assign n15185 = n15182 ^ n14738;
  assign n15186 = n15184 & n15185;
  assign n15187 = n15186 ^ n15182;
  assign n15188 = ~n14714 & ~n15187;
  assign n15189 = n15188 ^ n15182;
  assign n15181 = ~x6 & ~n14714;
  assign n15190 = n15189 ^ n15181;
  assign n15191 = n14737 ^ n14269;
  assign n15192 = n15191 ^ n15189;
  assign n15193 = n15189 ^ n15136;
  assign n15194 = n15189 & ~n15193;
  assign n15195 = n15194 ^ n15189;
  assign n15196 = n15192 & n15195;
  assign n15197 = n15196 ^ n15194;
  assign n15198 = n15197 ^ n15189;
  assign n15199 = n15198 ^ n15136;
  assign n15200 = ~n15190 & ~n15199;
  assign n15201 = n15200 ^ n15181;
  assign n15202 = n15201 ^ x7;
  assign n15203 = n15202 ^ n15179;
  assign n15204 = n15180 & ~n15203;
  assign n15205 = n15204 ^ n13862;
  assign n15206 = n15205 ^ n15154;
  assign n15207 = ~n15155 & n15206;
  assign n15208 = n15207 ^ n13444;
  assign n15209 = n15208 ^ n15151;
  assign n15210 = n15152 & ~n15209;
  assign n15211 = n15210 ^ n13031;
  assign n15212 = n15211 ^ n12617;
  assign n15213 = n14781 & ~n15136;
  assign n15214 = n15213 ^ n14784;
  assign n15215 = n15214 ^ n15211;
  assign n15216 = n15212 & n15215;
  assign n15217 = n15216 ^ n12617;
  assign n15218 = n15217 ^ n12230;
  assign n15219 = n14788 & ~n15136;
  assign n15220 = n15219 ^ n14790;
  assign n15221 = n15220 ^ n15217;
  assign n15222 = n15218 & ~n15221;
  assign n15223 = n15222 ^ n12230;
  assign n15224 = n15223 ^ n11820;
  assign n15225 = n14794 & ~n15136;
  assign n15226 = n15225 ^ n14796;
  assign n15227 = n15226 ^ n15223;
  assign n15228 = n15224 & n15227;
  assign n15229 = n15228 ^ n11820;
  assign n15230 = n15229 ^ n11395;
  assign n15231 = n14800 & ~n15136;
  assign n15232 = n15231 ^ n14802;
  assign n15233 = n15232 ^ n15229;
  assign n15234 = n15230 & ~n15233;
  assign n15235 = n15234 ^ n11395;
  assign n15236 = n15235 ^ n10956;
  assign n15237 = n14805 ^ n11395;
  assign n15238 = ~n15136 & n15237;
  assign n15239 = n15238 ^ n14735;
  assign n15240 = n15239 ^ n15235;
  assign n15241 = n15236 & n15240;
  assign n15242 = n15241 ^ n10956;
  assign n15243 = n15242 ^ n10585;
  assign n15244 = n14808 ^ n10956;
  assign n15245 = ~n15136 & n15244;
  assign n15246 = n15245 ^ n14731;
  assign n15247 = n15246 ^ n15242;
  assign n15248 = ~n15243 & ~n15247;
  assign n15249 = n15248 ^ n10585;
  assign n15250 = n15249 ^ n10229;
  assign n15251 = n14811 ^ n10585;
  assign n15252 = ~n15136 & ~n15251;
  assign n15253 = n15252 ^ n14727;
  assign n15254 = n15253 ^ n15249;
  assign n15255 = ~n15250 & ~n15254;
  assign n15256 = n15255 ^ n10229;
  assign n15257 = n15256 ^ n9867;
  assign n15258 = n14814 & ~n14823;
  assign n15259 = n15258 ^ n10229;
  assign n15260 = ~n15136 & ~n15259;
  assign n15261 = n15260 ^ n14817;
  assign n15262 = n15261 ^ n15256;
  assign n15263 = n15257 & ~n15262;
  assign n15264 = n15263 ^ n9867;
  assign n15265 = n15264 ^ n9502;
  assign n15266 = ~n14828 & ~n15136;
  assign n15267 = n15266 ^ n14830;
  assign n15268 = n15267 ^ n15264;
  assign n15269 = n15265 & ~n15268;
  assign n15270 = n15269 ^ n9502;
  assign n15271 = n15270 ^ n9129;
  assign n15272 = n14834 & ~n15136;
  assign n15273 = n15272 ^ n14836;
  assign n15274 = n15273 ^ n15270;
  assign n15275 = n15271 & ~n15274;
  assign n15276 = n15275 ^ n9129;
  assign n15277 = n15276 ^ n8769;
  assign n15278 = n14840 & ~n15136;
  assign n15279 = n15278 ^ n14843;
  assign n15280 = n15279 ^ n15276;
  assign n15281 = n15277 & n15280;
  assign n15282 = n15281 ^ n8769;
  assign n15283 = n15282 ^ n8422;
  assign n15284 = n14847 & ~n15136;
  assign n15285 = n15284 ^ n14849;
  assign n15286 = n15285 ^ n15282;
  assign n15287 = n15283 & ~n15286;
  assign n15288 = n15287 ^ n8422;
  assign n15289 = n15288 ^ n8083;
  assign n15290 = n14853 & ~n15136;
  assign n15291 = n15290 ^ n14855;
  assign n15292 = n15291 ^ n15288;
  assign n15293 = n15289 & n15292;
  assign n15294 = n15293 ^ n8083;
  assign n15295 = n15294 ^ n7777;
  assign n15296 = n14859 & ~n15136;
  assign n15297 = n15296 ^ n14861;
  assign n15298 = n15297 ^ n15294;
  assign n15299 = n15295 & ~n15298;
  assign n15300 = n15299 ^ n7777;
  assign n15301 = n15300 ^ n7463;
  assign n15302 = n14865 & ~n15136;
  assign n15303 = n15302 ^ n14867;
  assign n15304 = n15303 ^ n15300;
  assign n15305 = n15301 & n15304;
  assign n15306 = n15305 ^ n7463;
  assign n15307 = n15306 ^ n7135;
  assign n15308 = n14871 & ~n15136;
  assign n15309 = n15308 ^ n14873;
  assign n15310 = n15309 ^ n15306;
  assign n15311 = n15307 & ~n15310;
  assign n15312 = n15311 ^ n7135;
  assign n15313 = n15312 ^ n6802;
  assign n15314 = n14877 & ~n15136;
  assign n15315 = n15314 ^ n14879;
  assign n15316 = n15315 ^ n15312;
  assign n15317 = n15313 & ~n15316;
  assign n15318 = n15317 ^ n6802;
  assign n15319 = n15318 ^ n6479;
  assign n15320 = n14883 & ~n15136;
  assign n15321 = n15320 ^ n14885;
  assign n15322 = n15321 ^ n15318;
  assign n15323 = n15319 & ~n15322;
  assign n15324 = n15323 ^ n6479;
  assign n15325 = n15324 ^ n6181;
  assign n15326 = n14889 & ~n15136;
  assign n15327 = n15326 ^ n14891;
  assign n15328 = n15327 ^ n15324;
  assign n15329 = n15325 & n15328;
  assign n15330 = n15329 ^ n6181;
  assign n15331 = n15330 ^ n5905;
  assign n15332 = n14895 & ~n15136;
  assign n15333 = n15332 ^ n14897;
  assign n15334 = n15333 ^ n15330;
  assign n15335 = n15331 & ~n15334;
  assign n15336 = n15335 ^ n5905;
  assign n15337 = n15336 ^ n5625;
  assign n15338 = n14900 ^ n5905;
  assign n15339 = ~n15136 & n15338;
  assign n15340 = n15339 ^ n14724;
  assign n15341 = n15340 ^ n15336;
  assign n15342 = n15337 & n15341;
  assign n15343 = n15342 ^ n5625;
  assign n15344 = n15343 ^ n5363;
  assign n15345 = n14903 ^ n5625;
  assign n15346 = ~n15136 & n15345;
  assign n15347 = n15346 ^ n14716;
  assign n15348 = n15347 ^ n15343;
  assign n15349 = n15344 & ~n15348;
  assign n15350 = n15349 ^ n5363;
  assign n15351 = n15350 ^ n5108;
  assign n15352 = n14907 & ~n15136;
  assign n15353 = n15352 ^ n14909;
  assign n15354 = n15353 ^ n15350;
  assign n15355 = n15351 & n15354;
  assign n15356 = n15355 ^ n5108;
  assign n15357 = n15356 ^ n4851;
  assign n15358 = n14913 & ~n15136;
  assign n15359 = n15358 ^ n14915;
  assign n15360 = n15359 ^ n15356;
  assign n15361 = n15357 & ~n15360;
  assign n15362 = n15361 ^ n4851;
  assign n15363 = n15362 ^ n4606;
  assign n15364 = n14919 & ~n15136;
  assign n15365 = n15364 ^ n14921;
  assign n15366 = n15365 ^ n15362;
  assign n15367 = n15363 & n15366;
  assign n15368 = n15367 ^ n4606;
  assign n15369 = n15149 & n15368;
  assign n15370 = n15147 ^ n4133;
  assign n15371 = n4362 & n15144;
  assign n15372 = n15371 ^ n15147;
  assign n15373 = ~n15370 & n15372;
  assign n15374 = n15373 ^ n4133;
  assign n15375 = ~n15369 & ~n15374;
  assign n15376 = n15375 ^ n3882;
  assign n15377 = n14937 & ~n15136;
  assign n15378 = n15377 ^ n14939;
  assign n15379 = n15378 ^ n15375;
  assign n15380 = ~n15376 & n15379;
  assign n15381 = n15380 ^ n3882;
  assign n15382 = n15381 ^ n3634;
  assign n15383 = n14943 & ~n15136;
  assign n15384 = n15383 ^ n14945;
  assign n15385 = n15384 ^ n15381;
  assign n15386 = ~n15382 & n15385;
  assign n15387 = n15386 ^ n3634;
  assign n15388 = n15387 ^ n3397;
  assign n15389 = ~n14949 & ~n15136;
  assign n15390 = n15389 ^ n14951;
  assign n15391 = n15390 ^ n15387;
  assign n15392 = ~n15388 & n15391;
  assign n15393 = n15392 ^ n3397;
  assign n15394 = n15393 ^ n3177;
  assign n15395 = ~n14955 & ~n15136;
  assign n15396 = n15395 ^ n14957;
  assign n15397 = n15396 ^ n15393;
  assign n15398 = n15394 & n15397;
  assign n15399 = n15398 ^ n3177;
  assign n15400 = n15399 ^ n2980;
  assign n15401 = n14961 & ~n15136;
  assign n15402 = n15401 ^ n14963;
  assign n15403 = n15402 ^ n15399;
  assign n15404 = n15400 & ~n15403;
  assign n15405 = n15404 ^ n2980;
  assign n15406 = n15405 ^ n2782;
  assign n15407 = n14967 & ~n15136;
  assign n15408 = n15407 ^ n14969;
  assign n15409 = n15408 ^ n15405;
  assign n15410 = n15406 & ~n15409;
  assign n15411 = n15410 ^ n2782;
  assign n15412 = n15411 ^ n2583;
  assign n15413 = n14973 & ~n15136;
  assign n15414 = n15413 ^ n14975;
  assign n15415 = n15414 ^ n15411;
  assign n15416 = n15412 & ~n15415;
  assign n15417 = n15416 ^ n2583;
  assign n15418 = n15417 ^ n2374;
  assign n15419 = n14979 & ~n15136;
  assign n15420 = n15419 ^ n14981;
  assign n15421 = n15420 ^ n15417;
  assign n15422 = n15418 & n15421;
  assign n15423 = n15422 ^ n2374;
  assign n15424 = n15423 ^ n2194;
  assign n15425 = n14985 & ~n15136;
  assign n15426 = n15425 ^ n14987;
  assign n15427 = n15426 ^ n15423;
  assign n15428 = ~n15424 & ~n15427;
  assign n15429 = n15428 ^ n2194;
  assign n15430 = n15429 ^ n2011;
  assign n15431 = ~n14991 & ~n15136;
  assign n15432 = n15431 ^ n14993;
  assign n15433 = n15432 ^ n15429;
  assign n15434 = ~n15430 & ~n15433;
  assign n15435 = n15434 ^ n2011;
  assign n15436 = n15435 ^ n1804;
  assign n15437 = ~n14997 & ~n15136;
  assign n15438 = n15437 ^ n14999;
  assign n15439 = n15438 ^ n15435;
  assign n15440 = n15436 & ~n15439;
  assign n15441 = n15440 ^ n1804;
  assign n15442 = n15441 ^ n1621;
  assign n15443 = n15003 & ~n15136;
  assign n15444 = n15443 ^ n15005;
  assign n15445 = n15444 ^ n15441;
  assign n15446 = n15442 & n15445;
  assign n15447 = n15446 ^ n1621;
  assign n15448 = n15447 ^ n1458;
  assign n15449 = n15009 & ~n15136;
  assign n15450 = n15449 ^ n15011;
  assign n15451 = n15450 ^ n15447;
  assign n15452 = n15448 & ~n15451;
  assign n15453 = n15452 ^ n1458;
  assign n15454 = n15453 ^ n1299;
  assign n15455 = n15015 & ~n15136;
  assign n15456 = n15455 ^ n15017;
  assign n15457 = n15456 ^ n15453;
  assign n15458 = n15454 & n15457;
  assign n15459 = n15458 ^ n1299;
  assign n15460 = n15459 ^ n1158;
  assign n15461 = n15021 & ~n15136;
  assign n15462 = n15461 ^ n15024;
  assign n15463 = n15462 ^ n15459;
  assign n15464 = n15460 & ~n15463;
  assign n15465 = n15464 ^ n1158;
  assign n15466 = n15465 ^ n1027;
  assign n15467 = n15028 & ~n15136;
  assign n15468 = n15467 ^ n15031;
  assign n15469 = n15468 ^ n15465;
  assign n15470 = n15466 & n15469;
  assign n15471 = n15470 ^ n1027;
  assign n15472 = n15471 ^ n905;
  assign n15473 = n15035 & ~n15136;
  assign n15474 = n15473 ^ n15037;
  assign n15475 = n15474 ^ n15471;
  assign n15476 = n15472 & ~n15475;
  assign n15477 = n15476 ^ n905;
  assign n15478 = n15477 ^ n803;
  assign n15479 = n15041 & ~n15136;
  assign n15480 = n15479 ^ n15043;
  assign n15481 = n15480 ^ n15477;
  assign n15482 = n15478 & n15481;
  assign n15483 = n15482 ^ n803;
  assign n15484 = n15483 ^ n707;
  assign n15485 = n15047 & ~n15136;
  assign n15486 = n15485 ^ n15049;
  assign n15487 = n15486 ^ n15483;
  assign n15488 = ~n15484 & ~n15487;
  assign n15489 = n15488 ^ n707;
  assign n15490 = n15489 ^ n608;
  assign n15491 = ~n15053 & ~n15136;
  assign n15492 = n15491 ^ n15055;
  assign n15493 = n15492 ^ n15489;
  assign n15494 = ~n15490 & ~n15493;
  assign n15495 = n15494 ^ n608;
  assign n15496 = n15495 ^ n514;
  assign n15497 = ~n15059 & ~n15136;
  assign n15498 = n15497 ^ n15061;
  assign n15499 = n15498 ^ n15495;
  assign n15500 = n15496 & ~n15499;
  assign n15501 = n15500 ^ n514;
  assign n15502 = n15501 ^ n436;
  assign n15503 = n15065 & ~n15136;
  assign n15504 = n15503 ^ n15067;
  assign n15505 = n15504 ^ n15501;
  assign n15506 = n15502 & n15505;
  assign n15507 = n15506 ^ n436;
  assign n15508 = n15507 ^ n363;
  assign n15509 = n15071 & ~n15136;
  assign n15510 = n15509 ^ n15073;
  assign n15511 = n15510 ^ n15507;
  assign n15512 = n15508 & ~n15511;
  assign n15513 = n15512 ^ n363;
  assign n15514 = n15513 ^ n300;
  assign n15515 = n15077 & ~n15136;
  assign n15516 = n15515 ^ n15079;
  assign n15517 = n15516 ^ n15513;
  assign n15518 = n15514 & n15517;
  assign n15519 = n15518 ^ n300;
  assign n15520 = n15519 ^ n243;
  assign n15521 = n15083 & ~n15136;
  assign n15522 = n15521 ^ n15085;
  assign n15523 = n15522 ^ n15519;
  assign n15524 = n15520 & ~n15523;
  assign n15525 = n15524 ^ n243;
  assign n15526 = n15525 ^ n15141;
  assign n15527 = ~n15142 & n15526;
  assign n15528 = n15527 ^ n210;
  assign n15529 = n15528 ^ n15138;
  assign n15530 = ~n15139 & ~n15529;
  assign n15531 = n15530 ^ n147;
  assign n15532 = ~n132 & ~n15531;
  assign n15533 = ~n15119 & ~n15136;
  assign n15534 = n15533 ^ n15123;
  assign n15535 = ~n15532 & n15534;
  assign n15536 = n132 & n15531;
  assign n15538 = n15132 ^ n15097;
  assign n15539 = n15538 ^ n15097;
  assign n15540 = ~n14466 & ~n15107;
  assign n15541 = n15099 & ~n15540;
  assign n15542 = n15541 ^ n15097;
  assign n15543 = ~n15539 & ~n15542;
  assign n15544 = n15543 ^ n15097;
  assign n15545 = ~n133 & n15544;
  assign n15537 = ~n15535 & ~n15536;
  assign n15546 = n15545 ^ n15537;
  assign n15547 = n15127 & ~n15136;
  assign n15548 = n15547 ^ n15129;
  assign n15549 = n15548 ^ n15545;
  assign n15550 = n15549 ^ n15548;
  assign n15551 = ~n14466 & ~n14713;
  assign n15552 = n14701 & n15551;
  assign n15553 = n15099 & ~n15552;
  assign n15554 = ~n15538 & ~n15553;
  assign n15555 = n133 & ~n15554;
  assign n15556 = ~n15548 & n15555;
  assign n15557 = n15556 ^ n15548;
  assign n15558 = ~n15550 & n15557;
  assign n15559 = n15558 ^ n15548;
  assign n15560 = ~n15546 & ~n15559;
  assign n15561 = n15560 ^ n15537;
  assign n15562 = ~n15536 & n15561;
  assign n15563 = n15535 & n15562;
  assign n15564 = n15534 & ~n15548;
  assign n15565 = n15532 & ~n15564;
  assign n15566 = n133 & ~n15565;
  assign n15567 = ~n15563 & n15566;
  assign n15568 = n15536 ^ n15534;
  assign n15569 = n15561 & ~n15568;
  assign n15570 = ~n15548 & n15569;
  assign n15571 = n15570 ^ n15534;
  assign n15572 = n15567 & n15571;
  assign n15573 = n15548 ^ n15537;
  assign n15574 = n15561 ^ n15548;
  assign n15575 = n15561 ^ n133;
  assign n15576 = ~n15561 & n15575;
  assign n15577 = n15576 ^ n15561;
  assign n15578 = n15574 & ~n15577;
  assign n15579 = n15578 ^ n15576;
  assign n15580 = n15579 ^ n15561;
  assign n15581 = n15580 ^ n133;
  assign n15582 = n15573 & n15581;
  assign n15583 = n15582 ^ n133;
  assign n15584 = ~n15572 & n15583;
  assign n15585 = n15562 ^ n15534;
  assign n15586 = n15585 ^ n15534;
  assign n15587 = n15534 ^ n15532;
  assign n15588 = n15587 ^ n15534;
  assign n15589 = n15586 & ~n15588;
  assign n15590 = n15589 ^ n15534;
  assign n15591 = ~n133 & n15590;
  assign n15592 = n15525 ^ n210;
  assign n15593 = n15561 & n15592;
  assign n15594 = n15593 ^ n15141;
  assign n15595 = n15594 ^ n147;
  assign n15596 = n15520 & n15561;
  assign n15597 = n15596 ^ n15522;
  assign n15598 = n15597 ^ n210;
  assign n15599 = n15514 & n15561;
  assign n15600 = n15599 ^ n15516;
  assign n15601 = n15600 ^ n243;
  assign n15602 = n15508 & n15561;
  assign n15603 = n15602 ^ n15510;
  assign n15604 = n15603 ^ n300;
  assign n15605 = ~n15490 & n15561;
  assign n15606 = n15605 ^ n15492;
  assign n15607 = n514 & ~n15606;
  assign n15608 = n15496 & n15561;
  assign n15609 = n15608 ^ n15498;
  assign n15610 = n436 & n15609;
  assign n15611 = ~n15607 & ~n15610;
  assign n15612 = n15478 & n15561;
  assign n15613 = n15612 ^ n15480;
  assign n15614 = n15613 ^ n707;
  assign n15615 = n15472 & n15561;
  assign n15616 = n15615 ^ n15474;
  assign n15617 = n15616 ^ n803;
  assign n15618 = n15466 & n15561;
  assign n15619 = n15618 ^ n15468;
  assign n15620 = n15619 ^ n905;
  assign n15621 = n15460 & n15561;
  assign n15622 = n15621 ^ n15462;
  assign n15623 = n15622 ^ n1027;
  assign n15624 = n15454 & n15561;
  assign n15625 = n15624 ^ n15456;
  assign n15626 = n15625 ^ n1158;
  assign n15627 = n15448 & n15561;
  assign n15628 = n15627 ^ n15450;
  assign n15629 = n15628 ^ n1299;
  assign n15630 = n15442 & n15561;
  assign n15631 = n15630 ^ n15444;
  assign n15632 = n15631 ^ n1458;
  assign n15633 = n15436 & n15561;
  assign n15634 = n15633 ^ n15438;
  assign n15635 = n15634 ^ n1621;
  assign n15636 = ~n15430 & n15561;
  assign n15637 = n15636 ^ n15432;
  assign n15638 = n15637 ^ n1804;
  assign n15639 = n15418 & n15561;
  assign n15640 = n15639 ^ n15420;
  assign n15641 = n15640 ^ n2194;
  assign n15642 = n15412 & n15561;
  assign n15643 = n15642 ^ n15414;
  assign n15644 = n15643 ^ n2374;
  assign n15645 = n15400 & n15561;
  assign n15646 = n15645 ^ n15402;
  assign n15647 = n15646 ^ n2782;
  assign n15648 = n15394 & n15561;
  assign n15649 = n15648 ^ n15396;
  assign n15650 = n15649 ^ n2980;
  assign n15651 = ~n15388 & n15561;
  assign n15652 = n15651 ^ n15390;
  assign n15653 = n15652 ^ n3177;
  assign n15654 = ~n15382 & n15561;
  assign n15655 = n15654 ^ n15384;
  assign n15656 = n15655 ^ n3397;
  assign n15657 = ~n15376 & n15561;
  assign n15658 = n15657 ^ n15378;
  assign n15659 = n15658 ^ n3634;
  assign n15660 = n15368 ^ n4362;
  assign n15661 = n15561 & n15660;
  assign n15662 = n15661 ^ n15144;
  assign n15663 = n15662 ^ n4133;
  assign n15664 = n15363 & n15561;
  assign n15665 = n15664 ^ n15365;
  assign n15666 = n15665 ^ n4362;
  assign n15667 = n15351 & n15561;
  assign n15668 = n15667 ^ n15353;
  assign n15669 = n15668 ^ n4851;
  assign n15670 = n15337 & n15561;
  assign n15671 = n15670 ^ n15340;
  assign n15672 = n15671 ^ n5363;
  assign n15673 = n15331 & n15561;
  assign n15674 = n15673 ^ n15333;
  assign n15675 = n15674 ^ n5625;
  assign n15676 = n15325 & n15561;
  assign n15677 = n15676 ^ n15327;
  assign n15678 = n5905 & ~n15677;
  assign n15679 = n15678 ^ n15674;
  assign n15680 = n15675 & n15679;
  assign n15681 = n15680 ^ n15674;
  assign n15682 = n15681 ^ n15671;
  assign n15683 = n15682 ^ n15671;
  assign n15684 = n15236 & n15561;
  assign n15685 = n15684 ^ n15239;
  assign n15686 = ~n10585 & ~n15685;
  assign n15687 = n15230 & n15561;
  assign n15688 = n15687 ^ n15232;
  assign n15689 = n15688 ^ n10956;
  assign n15690 = n15224 & n15561;
  assign n15691 = n15690 ^ n15226;
  assign n15692 = n15691 ^ n11395;
  assign n15693 = n15218 & n15561;
  assign n15694 = n15693 ^ n15220;
  assign n15695 = n15694 ^ n11820;
  assign n15696 = n15212 & n15561;
  assign n15697 = n15696 ^ n15214;
  assign n15698 = n15697 ^ n12230;
  assign n15699 = n15208 ^ n13031;
  assign n15700 = n15561 & n15699;
  assign n15701 = n15700 ^ n15151;
  assign n15702 = n15701 ^ n12617;
  assign n15703 = n15205 ^ n13444;
  assign n15704 = n15561 & n15703;
  assign n15705 = n15704 ^ n15154;
  assign n15706 = n15705 ^ n13031;
  assign n15707 = n15180 & n15561;
  assign n15708 = n15707 ^ n15202;
  assign n15709 = n15708 ^ n13444;
  assign n15710 = n15176 ^ n14269;
  assign n15711 = n15561 & n15710;
  assign n15712 = n15711 ^ n15159;
  assign n15713 = n15712 ^ n13862;
  assign n15715 = n15169 ^ n15168;
  assign n15716 = n15715 ^ n15168;
  assign n15717 = n15168 ^ n15163;
  assign n15718 = n15717 ^ n15168;
  assign n15719 = n15716 & ~n15718;
  assign n15720 = n15719 ^ n15168;
  assign n15721 = n15136 & n15720;
  assign n15722 = n15721 ^ n15168;
  assign n15714 = ~x4 & ~n15136;
  assign n15723 = n15722 ^ n15714;
  assign n15724 = n15161 ^ n14714;
  assign n15725 = n15724 ^ n15722;
  assign n15726 = n15722 ^ n15561;
  assign n15727 = ~n15722 & ~n15726;
  assign n15728 = n15727 ^ n15722;
  assign n15729 = ~n15725 & ~n15728;
  assign n15730 = n15729 ^ n15727;
  assign n15731 = n15730 ^ n15722;
  assign n15732 = n15731 ^ n15561;
  assign n15733 = n15723 & ~n15732;
  assign n15734 = n15733 ^ n15714;
  assign n15735 = n15734 ^ x5;
  assign n15736 = n15735 ^ n14269;
  assign n15752 = n15161 ^ n15136;
  assign n15753 = n15561 & ~n15752;
  assign n15754 = n15753 ^ n15136;
  assign n15755 = n15754 ^ x4;
  assign n15737 = ~x0 & ~x1;
  assign n15738 = ~x2 & n15737;
  assign n15739 = n15136 & ~n15738;
  assign n15740 = n15561 ^ x3;
  assign n15741 = ~n15739 & ~n15740;
  assign n15742 = ~x3 & n15561;
  assign n15743 = n15742 ^ n15737;
  assign n15744 = n15743 ^ n15742;
  assign n15745 = n15742 ^ n15136;
  assign n15746 = n15745 ^ n15742;
  assign n15747 = n15744 & ~n15746;
  assign n15748 = n15747 ^ n15742;
  assign n15749 = ~x2 & n15748;
  assign n15750 = n15749 ^ n15742;
  assign n15751 = ~n15741 & ~n15750;
  assign n15756 = n15755 ^ n15751;
  assign n15757 = n15751 ^ n14714;
  assign n15758 = ~n15756 & n15757;
  assign n15759 = n15758 ^ n15751;
  assign n15760 = n15759 ^ n15735;
  assign n15761 = n15736 & n15760;
  assign n15762 = n15761 ^ n15735;
  assign n15763 = n15762 ^ n15712;
  assign n15764 = ~n15713 & ~n15763;
  assign n15765 = n15764 ^ n15712;
  assign n15766 = n15765 ^ n15708;
  assign n15767 = n15709 & ~n15766;
  assign n15768 = n15767 ^ n15708;
  assign n15769 = n15768 ^ n13031;
  assign n15770 = ~n15706 & n15769;
  assign n15771 = n15770 ^ n13031;
  assign n15772 = n15771 ^ n15701;
  assign n15773 = n15702 & n15772;
  assign n15774 = n15773 ^ n15701;
  assign n15775 = n15774 ^ n15697;
  assign n15776 = ~n15698 & ~n15775;
  assign n15777 = n15776 ^ n15697;
  assign n15778 = n15777 ^ n11820;
  assign n15779 = n15695 & ~n15778;
  assign n15780 = n15779 ^ n11820;
  assign n15781 = n15780 ^ n15691;
  assign n15782 = ~n15692 & n15781;
  assign n15783 = n15782 ^ n11395;
  assign n15784 = n15783 ^ n15688;
  assign n15785 = n15689 & ~n15784;
  assign n15786 = n15785 ^ n10956;
  assign n15787 = ~n15686 & ~n15786;
  assign n15788 = n10585 & n15685;
  assign n15789 = ~n15250 & n15561;
  assign n15790 = n15789 ^ n15253;
  assign n15791 = ~n9867 & n15790;
  assign n15792 = ~n15788 & ~n15791;
  assign n15793 = ~n15243 & n15561;
  assign n15794 = n15793 ^ n15246;
  assign n15795 = ~n10229 & ~n15794;
  assign n15796 = n15792 & ~n15795;
  assign n15797 = ~n15787 & n15796;
  assign n15798 = n15257 & n15561;
  assign n15799 = n15798 ^ n15261;
  assign n15800 = n9502 & n15799;
  assign n15801 = n15790 ^ n9867;
  assign n15802 = n10229 & n15794;
  assign n15803 = n15802 ^ n15790;
  assign n15804 = ~n15801 & ~n15803;
  assign n15805 = n15804 ^ n15790;
  assign n15806 = ~n15800 & n15805;
  assign n15807 = ~n15797 & n15806;
  assign n15808 = ~n9502 & ~n15799;
  assign n15809 = n15265 & n15561;
  assign n15810 = n15809 ^ n15267;
  assign n15811 = ~n9129 & ~n15810;
  assign n15812 = ~n15808 & ~n15811;
  assign n15813 = ~n15807 & n15812;
  assign n15814 = n9129 & n15810;
  assign n15815 = n15271 & n15561;
  assign n15816 = n15815 ^ n15273;
  assign n15817 = n8769 & n15816;
  assign n15818 = ~n15814 & ~n15817;
  assign n15819 = ~n15813 & n15818;
  assign n15820 = n15277 & n15561;
  assign n15821 = n15820 ^ n15279;
  assign n15822 = ~n8422 & n15821;
  assign n15823 = ~n8769 & ~n15816;
  assign n15824 = ~n15822 & ~n15823;
  assign n15825 = ~n15819 & n15824;
  assign n15826 = n8422 & ~n15821;
  assign n15827 = n15283 & n15561;
  assign n15828 = n15827 ^ n15285;
  assign n15829 = n8083 & n15828;
  assign n15830 = ~n15826 & ~n15829;
  assign n15831 = ~n15825 & n15830;
  assign n15832 = n15289 & n15561;
  assign n15833 = n15832 ^ n15291;
  assign n15834 = ~n7777 & n15833;
  assign n15835 = ~n8083 & ~n15828;
  assign n15836 = ~n15834 & ~n15835;
  assign n15837 = ~n15831 & n15836;
  assign n15838 = n7777 & ~n15833;
  assign n15839 = n15295 & n15561;
  assign n15840 = n15839 ^ n15297;
  assign n15841 = n7463 & n15840;
  assign n15842 = ~n15838 & ~n15841;
  assign n15843 = ~n15837 & n15842;
  assign n15844 = ~n7463 & ~n15840;
  assign n15845 = n15301 & n15561;
  assign n15846 = n15845 ^ n15303;
  assign n15847 = ~n7135 & n15846;
  assign n15848 = ~n15844 & ~n15847;
  assign n15849 = ~n15843 & n15848;
  assign n15850 = n7135 & ~n15846;
  assign n15851 = n15307 & n15561;
  assign n15852 = n15851 ^ n15309;
  assign n15853 = n6802 & n15852;
  assign n15854 = ~n15850 & ~n15853;
  assign n15855 = ~n15849 & n15854;
  assign n15856 = ~n6802 & ~n15852;
  assign n15857 = n15313 & n15561;
  assign n15858 = n15857 ^ n15315;
  assign n15859 = ~n6479 & ~n15858;
  assign n15860 = ~n15856 & ~n15859;
  assign n15861 = n15319 & n15561;
  assign n15862 = n15861 ^ n15321;
  assign n15863 = ~n6181 & ~n15862;
  assign n15864 = n15860 & ~n15863;
  assign n15865 = ~n15855 & n15864;
  assign n15866 = n15862 ^ n6181;
  assign n15867 = n6479 & n15858;
  assign n15868 = n15867 ^ n15862;
  assign n15869 = n15866 & ~n15868;
  assign n15870 = n15869 ^ n6181;
  assign n15871 = ~n15865 & ~n15870;
  assign n15872 = ~n5905 & n15677;
  assign n15873 = ~n5625 & ~n15674;
  assign n15874 = ~n15872 & ~n15873;
  assign n15875 = ~n15871 & n15874;
  assign n15876 = n15875 ^ n15671;
  assign n15877 = n15876 ^ n15671;
  assign n15878 = ~n15683 & ~n15877;
  assign n15879 = n15878 ^ n15671;
  assign n15880 = ~n15672 & ~n15879;
  assign n15881 = n15880 ^ n5363;
  assign n15882 = n15881 ^ n5108;
  assign n15883 = n15344 & n15561;
  assign n15884 = n15883 ^ n15347;
  assign n15885 = n15884 ^ n15881;
  assign n15886 = n15882 & n15885;
  assign n15887 = n15886 ^ n15881;
  assign n15888 = n15887 ^ n15668;
  assign n15889 = ~n15669 & n15888;
  assign n15890 = n15889 ^ n4851;
  assign n15891 = n15890 ^ n4606;
  assign n15892 = n15357 & n15561;
  assign n15893 = n15892 ^ n15359;
  assign n15894 = n15893 ^ n15890;
  assign n15895 = n15891 & n15894;
  assign n15896 = n15895 ^ n15890;
  assign n15897 = n15896 ^ n15665;
  assign n15898 = ~n15666 & n15897;
  assign n15899 = n15898 ^ n4362;
  assign n15900 = n15899 ^ n15662;
  assign n15901 = n15663 & ~n15900;
  assign n15902 = n15901 ^ n4133;
  assign n15903 = n15902 ^ n3882;
  assign n15904 = n15368 ^ n15144;
  assign n15905 = n15660 & ~n15904;
  assign n15906 = n15905 ^ n4362;
  assign n15907 = n15906 ^ n4133;
  assign n15908 = n15561 & n15907;
  assign n15909 = n15908 ^ n15147;
  assign n15910 = n15909 ^ n15902;
  assign n15911 = n15903 & ~n15910;
  assign n15912 = n15911 ^ n15902;
  assign n15913 = n15912 ^ n15658;
  assign n15914 = ~n15659 & n15913;
  assign n15915 = n15914 ^ n15658;
  assign n15916 = n15915 ^ n15655;
  assign n15917 = ~n15656 & ~n15916;
  assign n15918 = n15917 ^ n15655;
  assign n15919 = n15918 ^ n15652;
  assign n15920 = n15653 & ~n15919;
  assign n15921 = n15920 ^ n15652;
  assign n15922 = n15921 ^ n15649;
  assign n15923 = ~n15650 & n15922;
  assign n15924 = n15923 ^ n2980;
  assign n15925 = n15924 ^ n15646;
  assign n15926 = n15647 & ~n15925;
  assign n15927 = n15926 ^ n2782;
  assign n15928 = n15927 ^ n2583;
  assign n15929 = n15406 & n15561;
  assign n15930 = n15929 ^ n15408;
  assign n15931 = n15930 ^ n15927;
  assign n15932 = n15928 & n15931;
  assign n15933 = n15932 ^ n15927;
  assign n15934 = n15933 ^ n15643;
  assign n15935 = n15644 & ~n15934;
  assign n15936 = n15935 ^ n2374;
  assign n15937 = n15936 ^ n15640;
  assign n15938 = n15641 & n15937;
  assign n15939 = n15938 ^ n2194;
  assign n15940 = n15939 ^ n2011;
  assign n15941 = ~n15424 & n15561;
  assign n15942 = n15941 ^ n15426;
  assign n15943 = n15942 ^ n15939;
  assign n15944 = ~n15940 & ~n15943;
  assign n15945 = n15944 ^ n15939;
  assign n15946 = n15945 ^ n15637;
  assign n15947 = ~n15638 & n15946;
  assign n15948 = n15947 ^ n15637;
  assign n15949 = n15948 ^ n15634;
  assign n15950 = n15635 & ~n15949;
  assign n15951 = n15950 ^ n15634;
  assign n15952 = n15951 ^ n15631;
  assign n15953 = ~n15632 & ~n15952;
  assign n15954 = n15953 ^ n15631;
  assign n15955 = n15954 ^ n15628;
  assign n15956 = n15629 & ~n15955;
  assign n15957 = n15956 ^ n15628;
  assign n15958 = n15957 ^ n15625;
  assign n15959 = ~n15626 & ~n15958;
  assign n15960 = n15959 ^ n15625;
  assign n15961 = n15960 ^ n15622;
  assign n15962 = n15623 & ~n15961;
  assign n15963 = n15962 ^ n15622;
  assign n15964 = n15963 ^ n15619;
  assign n15965 = ~n15620 & ~n15964;
  assign n15966 = n15965 ^ n15619;
  assign n15967 = n15966 ^ n15616;
  assign n15968 = n15617 & n15967;
  assign n15969 = n15968 ^ n803;
  assign n15970 = n15969 ^ n15613;
  assign n15971 = n15614 & n15970;
  assign n15972 = n15971 ^ n707;
  assign n15973 = n15972 ^ n608;
  assign n15974 = ~n15484 & n15561;
  assign n15975 = n15974 ^ n15486;
  assign n15976 = n15975 ^ n15972;
  assign n15977 = ~n15973 & ~n15976;
  assign n15978 = n15977 ^ n15972;
  assign n15979 = n15611 & n15978;
  assign n15980 = n15609 ^ n436;
  assign n15981 = ~n514 & n15606;
  assign n15982 = n15981 ^ n15609;
  assign n15983 = n15980 & n15982;
  assign n15984 = n15983 ^ n436;
  assign n15985 = ~n15979 & n15984;
  assign n15986 = n15985 ^ n363;
  assign n15987 = n15502 & n15561;
  assign n15988 = n15987 ^ n15504;
  assign n15989 = n15988 ^ n15985;
  assign n15990 = n15986 & ~n15989;
  assign n15991 = n15990 ^ n15985;
  assign n15992 = n15991 ^ n15603;
  assign n15993 = n15604 & n15992;
  assign n15994 = n15993 ^ n15603;
  assign n15995 = n15994 ^ n15600;
  assign n15996 = ~n15601 & ~n15995;
  assign n15997 = n15996 ^ n15600;
  assign n15998 = n15997 ^ n15597;
  assign n15999 = n15598 & n15998;
  assign n16000 = n15999 ^ n210;
  assign n16001 = n16000 ^ n15594;
  assign n16002 = n15595 & n16001;
  assign n16003 = n16002 ^ n147;
  assign n16004 = n16003 ^ n132;
  assign n16005 = n15528 ^ n147;
  assign n16006 = n15561 & ~n16005;
  assign n16007 = n16006 ^ n15138;
  assign n16008 = n16007 ^ n16003;
  assign n16009 = n16004 & ~n16008;
  assign n16010 = n16009 ^ n16003;
  assign n16011 = ~n15591 & ~n16010;
  assign n16012 = ~n15584 & ~n16011;
  assign y0 = ~n16012;
  assign y1 = n15561;
  assign y2 = ~n15136;
  assign y3 = ~n14714;
  assign y4 = ~n14269;
  assign y5 = ~n13862;
  assign y6 = ~n13444;
  assign y7 = ~n13031;
  assign y8 = ~n12617;
  assign y9 = ~n12230;
  assign y10 = ~n11820;
  assign y11 = ~n11395;
  assign y12 = ~n10956;
  assign y13 = n10585;
  assign y14 = ~n10229;
  assign y15 = ~n9867;
  assign y16 = ~n9502;
  assign y17 = ~n9129;
  assign y18 = ~n8769;
  assign y19 = ~n8422;
  assign y20 = ~n8083;
  assign y21 = ~n7777;
  assign y22 = ~n7463;
  assign y23 = ~n7135;
  assign y24 = ~n6802;
  assign y25 = ~n6479;
  assign y26 = ~n6181;
  assign y27 = ~n5905;
  assign y28 = ~n5625;
  assign y29 = ~n5363;
  assign y30 = ~n5108;
  assign y31 = ~n4851;
  assign y32 = ~n4606;
  assign y33 = ~n4362;
  assign y34 = ~n4133;
  assign y35 = ~n3882;
  assign y36 = n3634;
  assign y37 = ~n3397;
  assign y38 = ~n3177;
  assign y39 = ~n2980;
  assign y40 = ~n2782;
  assign y41 = ~n2583;
  assign y42 = ~n2374;
  assign y43 = n2194;
  assign y44 = ~n2011;
  assign y45 = ~n1804;
  assign y46 = ~n1621;
  assign y47 = ~n1458;
  assign y48 = ~n1299;
  assign y49 = ~n1158;
  assign y50 = ~n1027;
  assign y51 = ~n905;
  assign y52 = ~n803;
  assign y53 = n707;
  assign y54 = ~n608;
  assign y55 = ~n514;
  assign y56 = ~n436;
  assign y57 = ~n363;
  assign y58 = ~n300;
  assign y59 = ~n243;
  assign y60 = ~n210;
  assign y61 = n147;
  assign y62 = n132;
  assign y63 = ~n133;
endmodule