module Xor(input logic a, b,
           output logic result);

    assign result = a ^ b;
    
endmodule