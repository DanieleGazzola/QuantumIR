module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701;
  assign n11 = ~x5 & ~x6;
  assign n20 = ~x0 & x7;
  assign n21 = ~x2 & ~x8;
  assign n22 = x2 & x8;
  assign n23 = ~x9 & n22;
  assign n24 = ~n21 & ~n23;
  assign n25 = n20 & ~n24;
  assign n26 = x0 & x9;
  assign n27 = ~x2 & x8;
  assign n28 = n26 & n27;
  assign n29 = ~n25 & ~n28;
  assign n30 = ~x3 & ~n29;
  assign n31 = x8 & x9;
  assign n32 = x2 & ~x3;
  assign n33 = n31 & n32;
  assign n34 = ~x8 & ~x9;
  assign n35 = ~x2 & x3;
  assign n36 = n34 & n35;
  assign n37 = ~n33 & ~n36;
  assign n38 = ~x0 & ~n37;
  assign n39 = x3 ^ x2;
  assign n40 = n39 ^ x0;
  assign n41 = x8 ^ x3;
  assign n42 = x9 ^ x3;
  assign n43 = n42 ^ x3;
  assign n44 = ~n41 & ~n43;
  assign n45 = n44 ^ x3;
  assign n46 = n45 ^ n39;
  assign n47 = ~n40 & n46;
  assign n48 = n47 ^ n44;
  assign n49 = n48 ^ x3;
  assign n50 = n49 ^ x0;
  assign n51 = ~n39 & ~n50;
  assign n52 = n51 ^ n39;
  assign n53 = ~n38 & n52;
  assign n54 = ~x7 & ~n53;
  assign n55 = ~n30 & ~n54;
  assign n56 = ~x1 & ~n55;
  assign n12 = ~x7 & ~x8;
  assign n13 = ~x2 & ~x3;
  assign n14 = ~x7 & ~x9;
  assign n15 = n13 & ~n14;
  assign n16 = ~x8 & x9;
  assign n17 = n16 ^ x0;
  assign n18 = n15 & n17;
  assign n19 = ~n12 & ~n18;
  assign n57 = n56 ^ n19;
  assign n58 = n11 & ~n57;
  assign n59 = ~x1 & ~x8;
  assign n60 = ~x3 & ~n59;
  assign n61 = ~x1 & n22;
  assign n62 = n61 ^ x8;
  assign n63 = x0 & ~n62;
  assign n64 = ~n60 & n63;
  assign n65 = ~x5 & ~x9;
  assign n66 = x8 ^ x2;
  assign n67 = n66 ^ n41;
  assign n68 = x8 ^ x1;
  assign n69 = n68 ^ n41;
  assign n70 = n41 & ~n69;
  assign n71 = n70 ^ n41;
  assign n72 = n67 & n71;
  assign n73 = n72 ^ n70;
  assign n74 = n73 ^ x8;
  assign n75 = n74 ^ n41;
  assign n76 = ~x0 & ~n75;
  assign n77 = n65 & ~n76;
  assign n78 = ~n64 & n77;
  assign n79 = ~x5 & x8;
  assign n80 = x0 & x1;
  assign n81 = x8 & n80;
  assign n82 = x8 ^ x5;
  assign n83 = n82 ^ x8;
  assign n84 = ~x1 & ~x2;
  assign n85 = n84 ^ x8;
  assign n86 = ~n83 & ~n85;
  assign n87 = n86 ^ x8;
  assign n88 = ~n13 & n87;
  assign n89 = ~n81 & ~n88;
  assign n90 = ~n79 & ~n89;
  assign n91 = n31 & ~n32;
  assign n92 = x5 & x9;
  assign n93 = ~n26 & ~n92;
  assign n94 = ~n91 & n93;
  assign n95 = ~x0 & ~x1;
  assign n96 = n35 ^ x8;
  assign n97 = ~n83 & n96;
  assign n98 = n97 ^ x8;
  assign n99 = n95 & n98;
  assign n100 = ~n94 & ~n99;
  assign n101 = ~n90 & n100;
  assign n102 = n13 & n95;
  assign n103 = x5 & n34;
  assign n104 = ~n102 & n103;
  assign n105 = x6 & ~x7;
  assign n106 = ~n104 & n105;
  assign n107 = ~n101 & n106;
  assign n108 = ~n78 & n107;
  assign n109 = ~x3 & ~n22;
  assign n110 = x0 & ~x1;
  assign n111 = ~x1 & x9;
  assign n112 = n111 ^ x2;
  assign n113 = n110 & n112;
  assign n114 = n109 & ~n113;
  assign n115 = x0 & ~x2;
  assign n116 = ~x9 & n115;
  assign n117 = x2 & n16;
  assign n118 = ~n116 & ~n117;
  assign n119 = x1 & ~n118;
  assign n120 = x3 & ~n27;
  assign n121 = ~n119 & n120;
  assign n122 = ~n114 & ~n121;
  assign n123 = x9 ^ x0;
  assign n124 = x1 & ~n123;
  assign n125 = x8 & ~n124;
  assign n126 = x5 & ~x6;
  assign n127 = ~x7 & n126;
  assign n128 = ~n125 & n127;
  assign n129 = ~n122 & n128;
  assign n130 = ~n108 & ~n129;
  assign n131 = ~n58 & n130;
  assign n133 = x6 ^ x5;
  assign n132 = n102 ^ x4;
  assign n134 = n133 ^ n132;
  assign n135 = n133 ^ n34;
  assign n136 = n133 & n135;
  assign n137 = n136 ^ n133;
  assign n138 = ~n134 & n137;
  assign n139 = n138 ^ n136;
  assign n140 = n139 ^ n133;
  assign n141 = n140 ^ n34;
  assign n142 = n102 & n141;
  assign n143 = n142 ^ n132;
  assign n144 = ~n131 & ~n143;
  assign n160 = n22 & n110;
  assign n161 = n21 & n95;
  assign n162 = n14 & ~n161;
  assign n163 = ~n160 & n162;
  assign n145 = ~x3 & ~x9;
  assign n146 = ~x0 & x8;
  assign n147 = x1 & ~x2;
  assign n148 = n146 & n147;
  assign n149 = ~x7 & x8;
  assign n150 = ~n21 & ~n149;
  assign n151 = n110 & ~n150;
  assign n152 = ~n148 & ~n151;
  assign n153 = n145 & ~n152;
  assign n154 = ~n95 & ~n115;
  assign n155 = ~x3 & ~n84;
  assign n156 = n31 ^ x7;
  assign n157 = n155 & n156;
  assign n158 = ~n154 & n157;
  assign n159 = ~n153 & ~n158;
  assign n164 = n163 ^ n159;
  assign n165 = n11 & ~n164;
  assign n166 = ~x1 & ~x5;
  assign n167 = x9 ^ x8;
  assign n168 = x3 ^ x0;
  assign n169 = n168 ^ x0;
  assign n170 = ~n123 & n169;
  assign n171 = n170 ^ x0;
  assign n172 = n167 & n171;
  assign n173 = n172 ^ x3;
  assign n174 = n166 & ~n173;
  assign n175 = x1 & ~n42;
  assign n176 = ~x9 & ~n79;
  assign n177 = n175 & ~n176;
  assign n178 = x2 & ~n92;
  assign n179 = ~n177 & n178;
  assign n180 = ~n174 & n179;
  assign n181 = n13 & n80;
  assign n182 = ~x2 & ~n65;
  assign n183 = ~n181 & ~n182;
  assign n184 = x1 & ~n146;
  assign n185 = n92 & n184;
  assign n186 = ~n183 & ~n185;
  assign n187 = ~x3 & ~n95;
  assign n188 = n16 & n80;
  assign n189 = n187 & ~n188;
  assign n190 = n16 & n110;
  assign n191 = x3 & ~n92;
  assign n192 = ~n190 & n191;
  assign n193 = ~n189 & ~n192;
  assign n194 = n186 & ~n193;
  assign n195 = n105 & ~n194;
  assign n196 = ~n180 & n195;
  assign n197 = ~x3 & n160;
  assign n198 = x2 & x3;
  assign n199 = n16 & n198;
  assign n200 = ~n145 & ~n199;
  assign n201 = x1 & ~n200;
  assign n202 = ~n197 & ~n201;
  assign n203 = ~n31 & ~n111;
  assign n204 = x9 & ~n13;
  assign n205 = n203 & ~n204;
  assign n206 = ~x0 & n205;
  assign n207 = x1 & ~n27;
  assign n208 = ~x9 & ~n32;
  assign n209 = ~n207 & n208;
  assign n210 = ~n206 & ~n209;
  assign n211 = n202 & n210;
  assign n212 = n127 & ~n211;
  assign n213 = ~n196 & ~n212;
  assign n214 = ~n165 & n213;
  assign n215 = ~x0 & ~x6;
  assign n216 = ~x9 & ~n215;
  assign n217 = ~x3 & n84;
  assign n218 = ~n216 & n217;
  assign n219 = n218 ^ n34;
  assign n220 = n219 ^ n218;
  assign n221 = n218 ^ n102;
  assign n222 = n221 ^ n218;
  assign n223 = ~n220 & n222;
  assign n224 = n223 ^ n218;
  assign n225 = ~x4 & ~n224;
  assign n226 = n225 ^ n218;
  assign n227 = ~n214 & n226;
  assign n264 = x1 & x9;
  assign n265 = x6 ^ x2;
  assign n266 = x8 ^ x6;
  assign n267 = n265 & n266;
  assign n268 = n267 ^ x2;
  assign n269 = n264 & ~n268;
  assign n270 = ~x0 & ~n269;
  assign n271 = ~x3 & x9;
  assign n272 = x0 & ~n21;
  assign n273 = n271 & ~n272;
  assign n258 = x1 & ~x6;
  assign n274 = x8 & ~x9;
  assign n275 = n258 & ~n274;
  assign n241 = x2 & ~x6;
  assign n276 = ~x3 & ~n241;
  assign n277 = ~n275 & n276;
  assign n278 = ~n273 & ~n277;
  assign n279 = ~n270 & ~n278;
  assign n280 = ~x7 & ~n279;
  assign n228 = x0 & ~n34;
  assign n229 = n147 & n228;
  assign n230 = ~x6 & x8;
  assign n231 = ~x1 & ~n230;
  assign n232 = n116 & n231;
  assign n233 = ~x0 & x2;
  assign n234 = n31 & n233;
  assign n235 = ~n232 & ~n234;
  assign n236 = ~n229 & n235;
  assign n237 = ~x2 & ~x6;
  assign n238 = ~x8 & ~n215;
  assign n239 = ~n237 & ~n238;
  assign n240 = x1 & ~x9;
  assign n242 = x0 & ~n241;
  assign n243 = n240 & ~n242;
  assign n244 = ~n239 & n243;
  assign n245 = ~x9 & ~n22;
  assign n246 = ~x6 & ~n31;
  assign n247 = n95 & ~n246;
  assign n248 = ~n245 & n247;
  assign n249 = ~n244 & ~n248;
  assign n250 = n236 & n249;
  assign n251 = ~x5 & ~x7;
  assign n252 = x0 & n240;
  assign n253 = n11 & ~n16;
  assign n254 = ~n252 & n253;
  assign n255 = ~n251 & ~n254;
  assign n256 = ~x3 & ~n20;
  assign n257 = ~n145 & ~n256;
  assign n259 = ~x0 & n14;
  assign n260 = n258 & n259;
  assign n261 = ~n257 & ~n260;
  assign n262 = ~n255 & n261;
  assign n263 = ~n250 & n262;
  assign n281 = n280 ^ n263;
  assign n287 = ~x1 & x8;
  assign n283 = ~x5 & x6;
  assign n288 = ~x6 & x9;
  assign n289 = ~n283 & ~n288;
  assign n290 = n287 & ~n289;
  assign n291 = ~n23 & n79;
  assign n292 = ~n146 & ~n291;
  assign n293 = ~n290 & n292;
  assign n294 = x2 & ~x5;
  assign n295 = ~n237 & ~n294;
  assign n296 = ~x1 & n295;
  assign n297 = n240 & n294;
  assign n298 = x5 & x6;
  assign n299 = ~x0 & ~n298;
  assign n300 = ~n182 & n299;
  assign n301 = ~n297 & n300;
  assign n302 = ~n296 & n301;
  assign n303 = ~n293 & ~n302;
  assign n304 = x1 & x6;
  assign n305 = n304 ^ x0;
  assign n306 = n304 ^ x9;
  assign n307 = n306 ^ x9;
  assign n308 = n294 ^ x9;
  assign n309 = n307 & n308;
  assign n310 = n309 ^ x9;
  assign n311 = n305 & n310;
  assign n312 = n295 ^ x0;
  assign n313 = n312 ^ x0;
  assign n314 = n313 ^ x8;
  assign n315 = x5 & n240;
  assign n316 = n315 ^ x9;
  assign n317 = ~x0 & n316;
  assign n318 = n317 ^ n315;
  assign n319 = n314 & ~n318;
  assign n320 = n319 ^ n317;
  assign n321 = n320 ^ n315;
  assign n322 = n321 ^ x0;
  assign n323 = ~x8 & n322;
  assign n324 = ~n311 & n323;
  assign n325 = ~n303 & ~n324;
  assign n282 = ~x2 & n95;
  assign n284 = ~x8 & n283;
  assign n285 = n282 & ~n284;
  assign n286 = n285 ^ x4;
  assign n326 = n325 ^ n286;
  assign n327 = n326 ^ n286;
  assign n328 = n286 ^ n285;
  assign n329 = ~n327 & ~n328;
  assign n330 = n329 ^ n286;
  assign n331 = x3 & ~n330;
  assign n332 = n331 ^ n286;
  assign n333 = n281 & ~n332;
  assign n334 = ~x0 & x5;
  assign n335 = ~n230 & n334;
  assign n336 = ~x5 & ~n274;
  assign n337 = x0 & ~n288;
  assign n338 = n336 & n337;
  assign n339 = ~n335 & ~n338;
  assign n340 = x1 & ~n339;
  assign n341 = x0 & x5;
  assign n342 = x1 & ~n341;
  assign n343 = ~x6 & n31;
  assign n344 = ~n342 & n343;
  assign n345 = n110 & ~n126;
  assign n346 = ~n336 & n345;
  assign n347 = ~n344 & ~n346;
  assign n348 = ~n340 & n347;
  assign n349 = ~n112 & ~n298;
  assign n350 = x3 & ~n349;
  assign n351 = ~n348 & n350;
  assign n352 = n34 ^ x2;
  assign n353 = n352 ^ n34;
  assign n354 = n167 ^ n34;
  assign n355 = ~n353 & n354;
  assign n356 = n355 ^ n34;
  assign n357 = x1 & n356;
  assign n358 = n84 ^ x1;
  assign n359 = n358 ^ x1;
  assign n360 = n34 ^ x1;
  assign n361 = n360 ^ x1;
  assign n362 = n359 & n361;
  assign n363 = n362 ^ x1;
  assign n364 = ~x6 & n363;
  assign n365 = n364 ^ x1;
  assign n366 = ~n357 & ~n365;
  assign n367 = n341 & ~n366;
  assign n368 = n31 & n95;
  assign n369 = ~x6 & ~n368;
  assign n370 = ~n241 & ~n369;
  assign n371 = n146 ^ x1;
  assign n372 = x9 ^ x1;
  assign n373 = n372 ^ n283;
  assign n374 = ~n371 & ~n373;
  assign n375 = n374 ^ n146;
  assign n376 = n283 & n375;
  assign n377 = n376 ^ x5;
  assign n378 = n370 & ~n377;
  assign n379 = n22 & n264;
  assign n380 = ~x6 & ~n379;
  assign n381 = ~n304 & n334;
  assign n382 = x2 & n283;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n380 & ~n383;
  assign n385 = ~n146 & n297;
  assign n386 = ~x3 & ~n385;
  assign n387 = ~n384 & n386;
  assign n388 = ~n378 & n387;
  assign n389 = ~n367 & n388;
  assign n390 = ~n133 & n217;
  assign n391 = n390 ^ x4;
  assign n392 = ~x7 & ~n391;
  assign n393 = ~n389 & n392;
  assign n394 = ~n351 & n393;
  assign n395 = ~x7 & n298;
  assign n396 = n95 ^ x2;
  assign n397 = n95 ^ x4;
  assign n398 = n397 ^ x4;
  assign n399 = n217 ^ x4;
  assign n400 = n399 ^ x4;
  assign n401 = n398 & n400;
  assign n402 = n401 ^ x4;
  assign n403 = n396 & ~n402;
  assign n404 = n395 & n403;
  assign n405 = x4 ^ x3;
  assign n406 = n282 ^ x4;
  assign n407 = n405 & ~n406;
  assign n408 = n395 & n407;
  assign n409 = ~x3 & ~x4;
  assign n471 = ~x2 & n251;
  assign n472 = ~n34 & n471;
  assign n473 = x6 & ~n472;
  assign n474 = x0 & ~n473;
  assign n475 = n379 ^ x5;
  assign n476 = n475 ^ n379;
  assign n477 = n476 ^ x7;
  assign n478 = n288 ^ x2;
  assign n479 = n288 & ~n478;
  assign n480 = n479 ^ n379;
  assign n481 = n480 ^ n288;
  assign n482 = n477 & ~n481;
  assign n483 = n482 ^ n479;
  assign n484 = n483 ^ n288;
  assign n485 = ~x7 & n484;
  assign n486 = n485 ^ x5;
  assign n487 = n474 & ~n486;
  assign n488 = ~x7 & ~n34;
  assign n489 = x2 & ~n488;
  assign n490 = n14 & n79;
  assign n491 = x7 & ~x8;
  assign n492 = x1 & ~n491;
  assign n493 = ~n490 & n492;
  assign n494 = ~n489 & n493;
  assign n495 = ~x2 & ~n14;
  assign n496 = ~n103 & ~n495;
  assign n497 = x7 & n31;
  assign n498 = ~x1 & ~n497;
  assign n499 = n496 & n498;
  assign n500 = ~n494 & ~n499;
  assign n501 = n487 & ~n500;
  assign n447 = n65 & ~n304;
  assign n448 = n149 & ~n447;
  assign n449 = x2 & ~n448;
  assign n450 = x5 & ~n258;
  assign n451 = ~n264 & ~n450;
  assign n452 = ~x7 & ~n451;
  assign n453 = ~x5 & ~n31;
  assign n454 = ~x1 & ~x6;
  assign n455 = ~n149 & n454;
  assign n456 = n453 & n455;
  assign n457 = ~n452 & ~n456;
  assign n458 = n449 & n457;
  assign n459 = n12 & n304;
  assign n460 = ~x2 & ~n395;
  assign n461 = ~n459 & n460;
  assign n462 = n11 ^ x7;
  assign n463 = ~x8 & ~n462;
  assign n464 = x1 & n11;
  assign n465 = n464 ^ x9;
  assign n466 = n463 & ~n465;
  assign n467 = n466 ^ n464;
  assign n468 = ~x9 & n467;
  assign n469 = n461 & ~n468;
  assign n470 = ~n458 & ~n469;
  assign n502 = n501 ^ n470;
  assign n410 = x4 & n102;
  assign n411 = x5 & ~x8;
  assign n412 = ~n80 & n411;
  assign n413 = ~n147 & n412;
  assign n414 = ~n116 & n413;
  assign n415 = n111 & n233;
  assign n416 = x5 & x8;
  assign n417 = ~n240 & n416;
  assign n418 = ~n415 & n417;
  assign n419 = ~x4 & ~n418;
  assign n420 = ~n414 & n419;
  assign n421 = n420 ^ x5;
  assign n422 = n420 ^ x6;
  assign n423 = n422 ^ x6;
  assign n424 = ~n22 & ~n288;
  assign n425 = x0 & ~n424;
  assign n426 = ~x1 & ~n16;
  assign n427 = ~x2 & x6;
  assign n428 = ~x0 & ~x9;
  assign n429 = n428 ^ n146;
  assign n430 = n427 & n429;
  assign n431 = n430 ^ n428;
  assign n432 = n426 & ~n431;
  assign n433 = ~n425 & n432;
  assign n434 = ~x0 & n31;
  assign n435 = ~n268 & n434;
  assign n436 = ~x2 & ~n146;
  assign n437 = n216 & n436;
  assign n438 = x1 & ~n437;
  assign n439 = ~n435 & n438;
  assign n440 = ~n433 & ~n439;
  assign n441 = n440 ^ x6;
  assign n442 = n423 & n441;
  assign n443 = n442 ^ x6;
  assign n444 = n421 & ~n443;
  assign n445 = n444 ^ x5;
  assign n446 = ~n410 & ~n445;
  assign n503 = n502 ^ n446;
  assign n504 = n503 ^ n502;
  assign n505 = n502 ^ x7;
  assign n506 = n505 ^ n502;
  assign n507 = ~n504 & ~n506;
  assign n508 = n507 ^ n502;
  assign n509 = ~n409 & n508;
  assign n510 = n509 ^ n502;
  assign n511 = ~n60 & ~n287;
  assign n512 = ~n203 & n511;
  assign n513 = x8 & n124;
  assign n514 = ~x3 & ~n513;
  assign n515 = ~n95 & ~n434;
  assign n516 = ~n514 & n515;
  assign n517 = ~n512 & n516;
  assign n518 = ~x2 & ~n517;
  assign n519 = n22 & n42;
  assign n520 = x0 & ~x8;
  assign n521 = ~n271 & n520;
  assign n522 = ~n35 & n521;
  assign n523 = ~n519 & ~n522;
  assign n524 = x1 & ~n523;
  assign n525 = n167 & n454;
  assign n526 = ~x0 & n13;
  assign n527 = n526 ^ x3;
  assign n528 = n525 & ~n527;
  assign n529 = n126 & ~n528;
  assign n530 = ~n524 & n529;
  assign n531 = ~n518 & n530;
  assign n582 = n34 & n187;
  assign n583 = n203 & ~n287;
  assign n584 = ~n582 & n583;
  assign n585 = ~n111 & n228;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~x2 & ~n586;
  assign n588 = x2 & ~n34;
  assign n589 = ~x0 & x3;
  assign n590 = ~n167 & n589;
  assign n591 = ~n588 & ~n590;
  assign n592 = ~x1 & ~n591;
  assign n593 = ~n33 & ~n592;
  assign n594 = ~n587 & n593;
  assign n533 = x2 ^ x0;
  assign n539 = x1 ^ x0;
  assign n540 = n539 ^ n42;
  assign n541 = n540 ^ x3;
  assign n532 = n42 ^ x1;
  assign n534 = n533 ^ n532;
  assign n542 = n541 ^ n534;
  assign n543 = n542 ^ n533;
  assign n544 = n533 & n543;
  assign n545 = n544 ^ n42;
  assign n546 = n545 ^ n534;
  assign n547 = n546 ^ n533;
  assign n548 = n547 ^ x3;
  assign n549 = n534 ^ n533;
  assign n550 = n549 ^ x3;
  assign n551 = n546 & n550;
  assign n552 = n551 ^ n42;
  assign n553 = n552 ^ n534;
  assign n554 = n553 ^ n533;
  assign n555 = n554 ^ x3;
  assign n556 = n548 & n555;
  assign n535 = n534 ^ n42;
  assign n536 = n535 ^ n533;
  assign n537 = n536 ^ x3;
  assign n538 = n536 & n537;
  assign n557 = n556 ^ n538;
  assign n558 = n557 ^ n544;
  assign n559 = n558 ^ n42;
  assign n560 = n559 ^ n534;
  assign n561 = n560 ^ n533;
  assign n562 = n561 ^ x3;
  assign n563 = x8 & n562;
  assign n564 = n41 ^ n39;
  assign n565 = n428 ^ x3;
  assign n566 = n565 ^ n41;
  assign n567 = n41 & ~n566;
  assign n568 = n567 ^ n41;
  assign n569 = n564 & n568;
  assign n570 = n569 ^ n567;
  assign n571 = n570 ^ x3;
  assign n572 = n571 ^ n41;
  assign n573 = n572 ^ x9;
  assign n574 = n573 ^ n572;
  assign n575 = n572 ^ n32;
  assign n576 = n575 ^ n572;
  assign n577 = n574 & n576;
  assign n578 = n577 ^ n572;
  assign n579 = x1 & ~n578;
  assign n580 = n579 ^ n572;
  assign n581 = ~n563 & n580;
  assign n595 = n594 ^ n581;
  assign n596 = n595 ^ n594;
  assign n597 = n594 ^ x6;
  assign n598 = n597 ^ n594;
  assign n599 = ~n596 & ~n598;
  assign n600 = n599 ^ n594;
  assign n601 = ~x4 & ~n600;
  assign n602 = n601 ^ x6;
  assign n603 = ~x5 & ~n602;
  assign n604 = ~n531 & ~n603;
  assign n605 = x4 & ~n102;
  assign n606 = x7 & ~n528;
  assign n607 = n14 & n27;
  assign n608 = ~n491 & ~n607;
  assign n609 = x0 & n454;
  assign n610 = ~n608 & n609;
  assign n611 = ~n606 & ~n610;
  assign n612 = ~n605 & n611;
  assign n613 = ~n604 & n612;
  assign n614 = n251 & n410;
  assign n615 = ~n11 & ~n246;
  assign n616 = ~n26 & ~n315;
  assign n617 = n539 ^ x8;
  assign n618 = n68 ^ x8;
  assign n619 = ~n167 & ~n618;
  assign n620 = n619 ^ x8;
  assign n621 = ~n617 & n620;
  assign n622 = n621 ^ x1;
  assign n623 = n616 & n622;
  assign n624 = ~x2 & ~n623;
  assign n625 = ~x1 & ~n245;
  assign n626 = ~n453 & n625;
  assign n627 = n386 & ~n626;
  assign n628 = ~n624 & n627;
  assign n629 = ~n615 & n628;
  assign n630 = ~n282 & ~n454;
  assign n631 = ~x9 & ~n238;
  assign n632 = ~n630 & n631;
  assign n633 = x9 & n265;
  assign n634 = ~n184 & n633;
  assign n635 = n237 & ~n287;
  assign n636 = x3 & ~x5;
  assign n637 = ~n635 & n636;
  assign n638 = ~n634 & n637;
  assign n639 = ~n632 & n638;
  assign n640 = n35 & n126;
  assign n641 = n583 ^ n95;
  assign n642 = n641 ^ n583;
  assign n643 = n583 ^ n31;
  assign n644 = n642 & n643;
  assign n645 = n644 ^ n583;
  assign n646 = n640 & ~n645;
  assign n647 = ~n639 & ~n646;
  assign n648 = ~n629 & n647;
  assign n649 = n11 & ~n31;
  assign n650 = ~x2 & ~n240;
  assign n651 = n95 & n588;
  assign n652 = ~n650 & ~n651;
  assign n653 = n649 & ~n652;
  assign n654 = x7 & ~n653;
  assign n655 = ~x4 & ~n654;
  assign n656 = ~n648 & n655;
  assign n657 = ~n614 & ~n656;
  assign n658 = ~n369 & n377;
  assign n659 = ~x1 & ~n34;
  assign n660 = n515 & ~n659;
  assign n661 = n11 & n660;
  assign n662 = ~n658 & ~n661;
  assign n663 = x5 ^ x2;
  assign n664 = n663 ^ x6;
  assign n665 = n298 & ~n664;
  assign n666 = n665 ^ n664;
  assign n667 = ~n662 & n666;
  assign n668 = x3 & ~x7;
  assign n669 = ~n667 & n668;
  assign n670 = n241 & n583;
  assign n671 = ~n11 & ~n84;
  assign n672 = ~n670 & n671;
  assign n673 = x7 ^ x2;
  assign n674 = n539 ^ x0;
  assign n675 = ~x9 & ~n146;
  assign n676 = n675 ^ x0;
  assign n677 = n674 & ~n676;
  assign n678 = n677 ^ x0;
  assign n679 = n678 ^ x7;
  assign n680 = n673 & ~n679;
  assign n681 = n680 ^ n677;
  assign n682 = n681 ^ x0;
  assign n683 = n682 ^ x2;
  assign n684 = ~x7 & ~n683;
  assign n685 = n684 ^ x7;
  assign n686 = n685 ^ x7;
  assign n687 = ~n651 & ~n686;
  assign n688 = n22 & n111;
  assign n689 = ~x3 & ~n688;
  assign n690 = ~n390 & n689;
  assign n691 = ~n687 & n690;
  assign n692 = ~n672 & n691;
  assign n693 = ~n669 & ~n692;
  assign n694 = ~n399 & ~n693;
  assign n695 = ~x7 & n11;
  assign n696 = n132 ^ n102;
  assign n697 = n198 & n660;
  assign n698 = n697 ^ n102;
  assign n699 = ~n696 & n698;
  assign n700 = n699 ^ n102;
  assign n701 = n695 & n700;
  assign y0 = n144;
  assign y1 = n227;
  assign y2 = n333;
  assign y3 = n394;
  assign y4 = n404;
  assign y5 = n408;
  assign y6 = ~n510;
  assign y7 = ~n613;
  assign y8 = n657;
  assign y9 = n694;
  assign y10 = n701;
endmodule