module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255, y256, y257, y258, y259, y260, y261, y262, y263, y264, y265, y266, y267, y268, y269, y270, y271, y272, y273, y274, y275, y276, y277, y278, y279, y280, y281, y282, y283, y284, y285, y286, y287, y288, y289, y290, y291, y292, y293, y294, y295, y296, y297, y298, y299, y300, y301, y302, y303, y304, y305, y306, y307, y308, y309, y310, y311, y312, y313, y314, y315, y316, y317, y318, y319, y320, y321, y322, y323, y324, y325, y326, y327, y328, y329, y330, y331, y332, y333, y334, y335, y336, y337, y338, y339, y340, y341, y342, y343, y344, y345, y346, y347, y348, y349, y350, y351, y352, y353, y354, y355, y356, y357, y358, y359, y360, y361, y362, y363, y364, y365, y366, y367, y368, y369, y370, y371, y372, y373, y374, y375, y376, y377, y378, y379, y380, y381, y382, y383, y384, y385, y386, y387, y388, y389, y390, y391, y392, y393, y394, y395, y396, y397, y398, y399, y400, y401, y402, y403, y404, y405, y406, y407, y408, y409, y410, y411, y412, y413, y414, y415, y416, y417, y418, y419, y420, y421, y422, y423, y424, y425, y426, y427, y428, y429, y430, y431, y432, y433, y434, y435, y436, y437, y438, y439, y440, y441, y442, y443, y444, y445, y446, y447, y448, y449, y450, y451, y452, y453, y454, y455, y456, y457, y458, y459, y460, y461, y462, y463, y464, y465, y466, y467, y468, y469, y470, y471, y472, y473, y474, y475, y476, y477, y478, y479, y480, y481, y482, y483, y484, y485, y486, y487, y488, y489, y490, y491, y492, y493, y494, y495, y496, y497, y498, y499, y500, y501, y502, y503, y504, y505, y506, y507, y508, y509, y510, y511, y512, y513, y514, y515, y516, y517, y518, y519, y520, y521, y522, y523, y524, y525, y526, y527, y528, y529, y530, y531, y532, y533, y534, y535, y536, y537, y538, y539, y540, y541, y542, y543, y544, y545, y546, y547, y548, y549, y550, y551, y552, y553, y554, y555, y556, y557, y558, y559, y560, y561, y562, y563, y564, y565, y566, y567, y568, y569, y570, y571, y572, y573, y574, y575, y576, y577, y578, y579, y580, y581, y582, y583, y584, y585, y586, y587, y588, y589, y590, y591, y592, y593, y594, y595, y596, y597, y598, y599, y600, y601, y602, y603, y604, y605, y606, y607, y608, y609, y610, y611, y612, y613, y614, y615, y616, y617, y618, y619, y620, y621, y622, y623, y624, y625, y626, y627, y628, y629, y630, y631, y632, y633, y634, y635, y636, y637, y638, y639, y640, y641, y642, y643, y644, y645, y646, y647, y648, y649, y650, y651, y652, y653, y654, y655, y656, y657, y658, y659, y660, y661, y662, y663, y664, y665, y666, y667, y668, y669, y670, y671, y672, y673, y674, y675, y676, y677, y678, y679, y680, y681, y682, y683, y684, y685, y686, y687, y688, y689, y690, y691, y692, y693, y694, y695, y696, y697, y698, y699, y700, y701, y702, y703, y704, y705, y706, y707, y708, y709, y710, y711, y712, y713, y714, y715, y716, y717, y718, y719, y720, y721, y722, y723, y724, y725, y726, y727, y728, y729, y730, y731, y732, y733, y734, y735, y736, y737, y738, y739, y740, y741, y742, y743, y744, y745, y746, y747, y748, y749, y750, y751, y752, y753, y754, y755, y756, y757, y758, y759, y760, y761, y762, y763, y764, y765, y766, y767, y768, y769, y770, y771, y772, y773, y774, y775, y776, y777, y778, y779, y780, y781, y782, y783, y784, y785, y786, y787, y788, y789, y790, y791, y792, y793, y794, y795, y796, y797, y798, y799, y800, y801, y802, y803, y804, y805, y806, y807, y808, y809, y810, y811, y812, y813, y814, y815, y816, y817, y818, y819, y820, y821, y822, y823, y824, y825, y826, y827, y828, y829, y830, y831, y832, y833, y834, y835, y836, y837, y838, y839, y840, y841, y842, y843, y844, y845, y846, y847, y848, y849, y850, y851, y852, y853, y854, y855, y856, y857, y858, y859, y860, y861, y862, y863, y864, y865, y866, y867, y868, y869, y870, y871, y872, y873, y874, y875, y876, y877, y878, y879, y880, y881, y882, y883, y884, y885, y886, y887, y888, y889, y890, y891, y892, y893, y894, y895, y896, y897, y898, y899, y900, y901, y902, y903, y904, y905, y906, y907, y908, y909, y910, y911, y912, y913, y914, y915, y916, y917, y918, y919, y920, y921, y922, y923, y924, y925, y926, y927, y928, y929, y930, y931, y932, y933, y934, y935, y936, y937, y938, y939, y940, y941, y942, y943, y944, y945, y946, y947, y948, y949, y950, y951, y952, y953, y954, y955, y956, y957, y958, y959, y960, y961, y962, y963, y964, y965, y966, y967, y968, y969, y970, y971, y972, y973, y974, y975, y976, y977, y978, y979, y980, y981, y982, y983, y984, y985, y986, y987, y988, y989, y990, y991, y992, y993, y994, y995, y996, y997, y998, y999, y1000, y1001, y1002, y1003, y1004, y1005, y1006, y1007, y1008, y1009, y1010, y1011, y1012, y1013, y1014, y1015, y1016, y1017, y1018, y1019, y1020, y1021, y1022, y1023, y1024, y1025, y1026, y1027, y1028, y1029, y1030, y1031, y1032, y1033, y1034, y1035, y1036, y1037, y1038, y1039, y1040, y1041, y1042, y1043, y1044, y1045, y1046, y1047, y1048, y1049, y1050, y1051, y1052, y1053, y1054, y1055, y1056, y1057, y1058, y1059, y1060, y1061, y1062, y1063, y1064, y1065, y1066, y1067, y1068, y1069, y1070, y1071, y1072, y1073, y1074, y1075, y1076, y1077, y1078, y1079, y1080, y1081, y1082, y1083, y1084, y1085, y1086, y1087, y1088, y1089, y1090, y1091, y1092, y1093, y1094, y1095, y1096, y1097, y1098, y1099, y1100, y1101, y1102, y1103, y1104, y1105, y1106, y1107, y1108, y1109, y1110, y1111, y1112, y1113, y1114, y1115, y1116, y1117, y1118, y1119, y1120, y1121, y1122, y1123, y1124, y1125, y1126, y1127, y1128, y1129, y1130, y1131, y1132, y1133, y1134, y1135, y1136, y1137, y1138, y1139, y1140, y1141, y1142, y1143, y1144, y1145, y1146, y1147, y1148, y1149, y1150, y1151, y1152, y1153, y1154, y1155, y1156, y1157, y1158, y1159, y1160, y1161, y1162, y1163, y1164, y1165, y1166, y1167, y1168, y1169, y1170, y1171, y1172, y1173, y1174, y1175, y1176, y1177, y1178, y1179, y1180, y1181, y1182, y1183, y1184, y1185, y1186, y1187, y1188, y1189, y1190, y1191, y1192, y1193, y1194, y1195, y1196, y1197, y1198, y1199, y1200, y1201, y1202, y1203, y1204, y1205, y1206, y1207, y1208, y1209, y1210, y1211, y1212, y1213, y1214, y1215, y1216, y1217, y1218, y1219, y1220, y1221, y1222, y1223, y1224, y1225, y1226, y1227, y1228, y1229, y1230);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255, y256, y257, y258, y259, y260, y261, y262, y263, y264, y265, y266, y267, y268, y269, y270, y271, y272, y273, y274, y275, y276, y277, y278, y279, y280, y281, y282, y283, y284, y285, y286, y287, y288, y289, y290, y291, y292, y293, y294, y295, y296, y297, y298, y299, y300, y301, y302, y303, y304, y305, y306, y307, y308, y309, y310, y311, y312, y313, y314, y315, y316, y317, y318, y319, y320, y321, y322, y323, y324, y325, y326, y327, y328, y329, y330, y331, y332, y333, y334, y335, y336, y337, y338, y339, y340, y341, y342, y343, y344, y345, y346, y347, y348, y349, y350, y351, y352, y353, y354, y355, y356, y357, y358, y359, y360, y361, y362, y363, y364, y365, y366, y367, y368, y369, y370, y371, y372, y373, y374, y375, y376, y377, y378, y379, y380, y381, y382, y383, y384, y385, y386, y387, y388, y389, y390, y391, y392, y393, y394, y395, y396, y397, y398, y399, y400, y401, y402, y403, y404, y405, y406, y407, y408, y409, y410, y411, y412, y413, y414, y415, y416, y417, y418, y419, y420, y421, y422, y423, y424, y425, y426, y427, y428, y429, y430, y431, y432, y433, y434, y435, y436, y437, y438, y439, y440, y441, y442, y443, y444, y445, y446, y447, y448, y449, y450, y451, y452, y453, y454, y455, y456, y457, y458, y459, y460, y461, y462, y463, y464, y465, y466, y467, y468, y469, y470, y471, y472, y473, y474, y475, y476, y477, y478, y479, y480, y481, y482, y483, y484, y485, y486, y487, y488, y489, y490, y491, y492, y493, y494, y495, y496, y497, y498, y499, y500, y501, y502, y503, y504, y505, y506, y507, y508, y509, y510, y511, y512, y513, y514, y515, y516, y517, y518, y519, y520, y521, y522, y523, y524, y525, y526, y527, y528, y529, y530, y531, y532, y533, y534, y535, y536, y537, y538, y539, y540, y541, y542, y543, y544, y545, y546, y547, y548, y549, y550, y551, y552, y553, y554, y555, y556, y557, y558, y559, y560, y561, y562, y563, y564, y565, y566, y567, y568, y569, y570, y571, y572, y573, y574, y575, y576, y577, y578, y579, y580, y581, y582, y583, y584, y585, y586, y587, y588, y589, y590, y591, y592, y593, y594, y595, y596, y597, y598, y599, y600, y601, y602, y603, y604, y605, y606, y607, y608, y609, y610, y611, y612, y613, y614, y615, y616, y617, y618, y619, y620, y621, y622, y623, y624, y625, y626, y627, y628, y629, y630, y631, y632, y633, y634, y635, y636, y637, y638, y639, y640, y641, y642, y643, y644, y645, y646, y647, y648, y649, y650, y651, y652, y653, y654, y655, y656, y657, y658, y659, y660, y661, y662, y663, y664, y665, y666, y667, y668, y669, y670, y671, y672, y673, y674, y675, y676, y677, y678, y679, y680, y681, y682, y683, y684, y685, y686, y687, y688, y689, y690, y691, y692, y693, y694, y695, y696, y697, y698, y699, y700, y701, y702, y703, y704, y705, y706, y707, y708, y709, y710, y711, y712, y713, y714, y715, y716, y717, y718, y719, y720, y721, y722, y723, y724, y725, y726, y727, y728, y729, y730, y731, y732, y733, y734, y735, y736, y737, y738, y739, y740, y741, y742, y743, y744, y745, y746, y747, y748, y749, y750, y751, y752, y753, y754, y755, y756, y757, y758, y759, y760, y761, y762, y763, y764, y765, y766, y767, y768, y769, y770, y771, y772, y773, y774, y775, y776, y777, y778, y779, y780, y781, y782, y783, y784, y785, y786, y787, y788, y789, y790, y791, y792, y793, y794, y795, y796, y797, y798, y799, y800, y801, y802, y803, y804, y805, y806, y807, y808, y809, y810, y811, y812, y813, y814, y815, y816, y817, y818, y819, y820, y821, y822, y823, y824, y825, y826, y827, y828, y829, y830, y831, y832, y833, y834, y835, y836, y837, y838, y839, y840, y841, y842, y843, y844, y845, y846, y847, y848, y849, y850, y851, y852, y853, y854, y855, y856, y857, y858, y859, y860, y861, y862, y863, y864, y865, y866, y867, y868, y869, y870, y871, y872, y873, y874, y875, y876, y877, y878, y879, y880, y881, y882, y883, y884, y885, y886, y887, y888, y889, y890, y891, y892, y893, y894, y895, y896, y897, y898, y899, y900, y901, y902, y903, y904, y905, y906, y907, y908, y909, y910, y911, y912, y913, y914, y915, y916, y917, y918, y919, y920, y921, y922, y923, y924, y925, y926, y927, y928, y929, y930, y931, y932, y933, y934, y935, y936, y937, y938, y939, y940, y941, y942, y943, y944, y945, y946, y947, y948, y949, y950, y951, y952, y953, y954, y955, y956, y957, y958, y959, y960, y961, y962, y963, y964, y965, y966, y967, y968, y969, y970, y971, y972, y973, y974, y975, y976, y977, y978, y979, y980, y981, y982, y983, y984, y985, y986, y987, y988, y989, y990, y991, y992, y993, y994, y995, y996, y997, y998, y999, y1000, y1001, y1002, y1003, y1004, y1005, y1006, y1007, y1008, y1009, y1010, y1011, y1012, y1013, y1014, y1015, y1016, y1017, y1018, y1019, y1020, y1021, y1022, y1023, y1024, y1025, y1026, y1027, y1028, y1029, y1030, y1031, y1032, y1033, y1034, y1035, y1036, y1037, y1038, y1039, y1040, y1041, y1042, y1043, y1044, y1045, y1046, y1047, y1048, y1049, y1050, y1051, y1052, y1053, y1054, y1055, y1056, y1057, y1058, y1059, y1060, y1061, y1062, y1063, y1064, y1065, y1066, y1067, y1068, y1069, y1070, y1071, y1072, y1073, y1074, y1075, y1076, y1077, y1078, y1079, y1080, y1081, y1082, y1083, y1084, y1085, y1086, y1087, y1088, y1089, y1090, y1091, y1092, y1093, y1094, y1095, y1096, y1097, y1098, y1099, y1100, y1101, y1102, y1103, y1104, y1105, y1106, y1107, y1108, y1109, y1110, y1111, y1112, y1113, y1114, y1115, y1116, y1117, y1118, y1119, y1120, y1121, y1122, y1123, y1124, y1125, y1126, y1127, y1128, y1129, y1130, y1131, y1132, y1133, y1134, y1135, y1136, y1137, y1138, y1139, y1140, y1141, y1142, y1143, y1144, y1145, y1146, y1147, y1148, y1149, y1150, y1151, y1152, y1153, y1154, y1155, y1156, y1157, y1158, y1159, y1160, y1161, y1162, y1163, y1164, y1165, y1166, y1167, y1168, y1169, y1170, y1171, y1172, y1173, y1174, y1175, y1176, y1177, y1178, y1179, y1180, y1181, y1182, y1183, y1184, y1185, y1186, y1187, y1188, y1189, y1190, y1191, y1192, y1193, y1194, y1195, y1196, y1197, y1198, y1199, y1200, y1201, y1202, y1203, y1204, y1205, y1206, y1207, y1208, y1209, y1210, y1211, y1212, y1213, y1214, y1215, y1216, y1217, y1218, y1219, y1220, y1221, y1222, y1223, y1224, y1225, y1226, y1227, y1228, y1229, y1230;
  wire n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485;
  assign n1205 = x32 & ~x95;
  assign n1206 = ~x85 & ~x106;
  assign n1207 = ~x76 & n1206;
  assign n1208 = ~x48 & ~x61;
  assign n1209 = n1207 & n1208;
  assign n1210 = ~x104 & n1209;
  assign n1211 = ~x89 & n1210;
  assign n1212 = ~x49 & n1211;
  assign n1213 = ~x45 & n1212;
  assign n1214 = ~x69 & ~x83;
  assign n1215 = ~x103 & n1214;
  assign n1216 = ~x82 & ~x111;
  assign n1217 = ~x36 & n1216;
  assign n1218 = ~x66 & n1217;
  assign n1219 = n1215 & n1218;
  assign n1220 = n1213 & n1219;
  assign n1221 = ~x73 & n1220;
  assign n1222 = ~x88 & ~x98;
  assign n1223 = ~x102 & ~x107;
  assign n1224 = n1222 & n1223;
  assign n1225 = ~x64 & ~x65;
  assign n1226 = ~x63 & n1225;
  assign n1227 = n1224 & n1226;
  assign n1228 = ~x81 & n1227;
  assign n1229 = n1221 & n1228;
  assign n1230 = ~x67 & ~x68;
  assign n1231 = ~x71 & ~x84;
  assign n1232 = n1230 & n1231;
  assign n1233 = n1229 & n1232;
  assign n1234 = ~x91 & ~x109;
  assign n1235 = ~x46 & ~x47;
  assign n1236 = n1234 & n1235;
  assign n1237 = ~x77 & ~x86;
  assign n1238 = ~x50 & ~x110;
  assign n1239 = n1237 & n1238;
  assign n1240 = n1236 & n1239;
  assign n1241 = ~x53 & ~x60;
  assign n1242 = ~x58 & n1241;
  assign n1243 = ~x97 & ~x108;
  assign n1244 = ~x94 & n1243;
  assign n1245 = n1242 & n1244;
  assign n1246 = n1240 & n1245;
  assign n1247 = n1233 & n1246;
  assign n1248 = ~x72 & ~x96;
  assign n1249 = ~x51 & ~x70;
  assign n1250 = n1248 & n1249;
  assign n1251 = ~x35 & ~x93;
  assign n1252 = ~x90 & n1251;
  assign n1253 = n1250 & n1252;
  assign n1254 = n1247 & n1253;
  assign n1255 = ~x40 & n1254;
  assign n1256 = n1205 & n1255;
  assign n1257 = x210 ^ x198;
  assign n1258 = x299 & n1257;
  assign n1259 = n1258 ^ x198;
  assign n1260 = ~x841 & ~n1259;
  assign n1261 = x225 & ~n1260;
  assign n1262 = n1256 & n1261;
  assign n1263 = n1247 & n1252;
  assign n1264 = ~x32 & ~x95;
  assign n1265 = ~x40 & n1264;
  assign n1269 = x96 ^ x51;
  assign n1270 = x96 ^ x72;
  assign n1271 = n1270 ^ x70;
  assign n1272 = ~n1269 & n1271;
  assign n1274 = n1272 ^ n1265;
  assign n1266 = x72 ^ x70;
  assign n1267 = n1266 ^ x70;
  assign n1268 = ~n1266 & ~n1267;
  assign n1275 = n1268 ^ n1266;
  assign n1276 = ~n1274 & ~n1275;
  assign n1273 = n1272 ^ n1268;
  assign n1277 = n1276 ^ n1273;
  assign n1278 = ~n1265 & n1277;
  assign n1279 = n1278 ^ n1272;
  assign n1280 = n1279 ^ n1268;
  assign n1281 = n1280 ^ n1276;
  assign n1282 = n1263 & n1281;
  assign n1283 = x96 & n1282;
  assign n1284 = x95 & ~x479;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = n1250 & n1265;
  assign n1456 = x40 ^ x32;
  assign n1457 = n1456 ^ x95;
  assign n1458 = x40 & x95;
  assign n1459 = n1457 & n1458;
  assign n1460 = n1459 ^ n1457;
  assign n1287 = ~x50 & n1241;
  assign n1288 = ~x77 & n1287;
  assign n1289 = n1243 & n1288;
  assign n1290 = ~x86 & ~x94;
  assign n1291 = n1289 & n1290;
  assign n1292 = n1233 & n1291;
  assign n1293 = ~x46 & ~x109;
  assign n1294 = n1241 ^ x50;
  assign n1295 = x53 & x60;
  assign n1296 = ~x77 & ~n1295;
  assign n1297 = n1296 ^ n1241;
  assign n1298 = ~n1294 & n1297;
  assign n1299 = n1298 ^ n1241;
  assign n1300 = n1293 & n1299;
  assign n1301 = n1292 & n1300;
  assign n1302 = ~x58 & ~x90;
  assign n1303 = ~x47 & ~x110;
  assign n1304 = n1302 & n1303;
  assign n1305 = ~x91 & ~x93;
  assign n1306 = n1304 & n1305;
  assign n1307 = ~n1301 & ~n1306;
  assign n1308 = x91 ^ x47;
  assign n1309 = ~n1302 & n1308;
  assign n1310 = n1251 & ~n1309;
  assign n1311 = x91 & ~n1303;
  assign n1312 = n1310 & ~n1311;
  assign n1313 = x110 ^ x90;
  assign n1314 = x110 ^ x47;
  assign n1315 = x90 ^ x58;
  assign n1316 = n1315 ^ x110;
  assign n1317 = x110 & ~n1316;
  assign n1318 = n1317 ^ x110;
  assign n1319 = n1314 & n1318;
  assign n1320 = n1319 ^ n1317;
  assign n1321 = n1320 ^ x110;
  assign n1322 = n1321 ^ n1315;
  assign n1323 = n1313 & ~n1322;
  assign n1324 = n1323 ^ x110;
  assign n1325 = n1312 & ~n1324;
  assign n1326 = ~n1307 & n1325;
  assign n1327 = ~x46 & ~n1234;
  assign n1328 = n1327 ^ n1292;
  assign n1329 = n1328 ^ n1327;
  assign n1330 = ~x73 & ~x84;
  assign n1331 = ~x68 & n1330;
  assign n1332 = ~x66 & n1331;
  assign n1333 = n1213 & n1332;
  assign n1334 = n1215 & n1333;
  assign n1336 = x111 ^ x82;
  assign n1337 = n1336 ^ x36;
  assign n1335 = x67 ^ x36;
  assign n1338 = n1337 ^ n1335;
  assign n1339 = x82 ^ x67;
  assign n1340 = n1339 ^ x36;
  assign n1341 = n1340 ^ x36;
  assign n1342 = ~n1336 & n1341;
  assign n1343 = n1342 ^ n1336;
  assign n1344 = n1340 & ~n1343;
  assign n1345 = n1344 ^ x36;
  assign n1346 = n1338 & n1345;
  assign n1347 = n1346 ^ n1342;
  assign n1348 = n1347 ^ x36;
  assign n1349 = n1348 ^ n1335;
  assign n1350 = n1334 & ~n1349;
  assign n1351 = ~x36 & ~x67;
  assign n1352 = n1216 & n1351;
  assign n1353 = n1215 & n1352;
  assign n1354 = ~n1350 & ~n1353;
  assign n1355 = x104 & ~n1209;
  assign n1356 = ~x49 & ~n1355;
  assign n1357 = n1356 ^ x89;
  assign n1358 = n1210 ^ x89;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = n1359 ^ x89;
  assign n1361 = ~x45 & ~n1360;
  assign n1362 = ~n1212 & ~n1361;
  assign n1363 = x61 ^ x48;
  assign n1364 = n1207 & n1363;
  assign n1365 = x106 ^ x85;
  assign n1366 = x85 ^ x76;
  assign n1367 = n1365 & n1366;
  assign n1368 = n1367 ^ x85;
  assign n1369 = n1208 & ~n1368;
  assign n1370 = ~n1364 & ~n1369;
  assign n1371 = n1332 & ~n1370;
  assign n1372 = ~n1362 & n1371;
  assign n1373 = x68 ^ x66;
  assign n1374 = n1373 ^ x73;
  assign n1375 = n1374 ^ x84;
  assign n1376 = x73 ^ x68;
  assign n1377 = x84 ^ x68;
  assign n1378 = n1376 & n1377;
  assign n1379 = n1378 ^ x68;
  assign n1380 = n1375 & ~n1379;
  assign n1381 = n1213 & n1380;
  assign n1382 = ~n1372 & ~n1381;
  assign n1383 = ~n1354 & ~n1382;
  assign n1384 = n1333 & n1352;
  assign n1385 = x83 ^ x69;
  assign n1386 = x103 ^ x83;
  assign n1387 = n1385 & ~n1386;
  assign n1388 = n1387 ^ x69;
  assign n1389 = n1384 & ~n1388;
  assign n1390 = ~n1383 & ~n1389;
  assign n1391 = n1229 & n1384;
  assign n1392 = ~x71 & ~x81;
  assign n1393 = n1227 & n1392;
  assign n1394 = ~n1391 & ~n1393;
  assign n1395 = ~n1390 & ~n1394;
  assign n1396 = n1221 & n1232;
  assign n1401 = x98 ^ x88;
  assign n1402 = n1401 ^ x102;
  assign n1403 = n1402 ^ x107;
  assign n1404 = x107 ^ x98;
  assign n1405 = x102 ^ x98;
  assign n1406 = n1404 & n1405;
  assign n1407 = n1406 ^ x98;
  assign n1408 = n1403 & ~n1407;
  assign n1409 = n1408 ^ n1224;
  assign n1410 = ~x81 & n1409;
  assign n1411 = n1410 ^ n1224;
  assign n1397 = ~x102 & n1232;
  assign n1398 = ~x81 & n1222;
  assign n1399 = n1397 & n1398;
  assign n1412 = n1411 ^ n1399;
  assign n1413 = n1412 ^ x64;
  assign n1414 = n1413 ^ x63;
  assign n1415 = n1414 ^ x65;
  assign n1400 = n1399 ^ x65;
  assign n1416 = n1415 ^ n1400;
  assign n1418 = x64 ^ x63;
  assign n1419 = n1418 ^ n1415;
  assign n1417 = n1414 ^ x63;
  assign n1420 = n1419 ^ n1417;
  assign n1421 = n1416 & n1420;
  assign n1422 = n1421 ^ n1414;
  assign n1423 = n1422 ^ n1418;
  assign n1424 = n1423 ^ n1417;
  assign n1425 = n1419 ^ n1400;
  assign n1426 = n1422 & n1425;
  assign n1427 = n1426 ^ n1414;
  assign n1428 = n1427 ^ n1415;
  assign n1429 = n1428 ^ n1400;
  assign n1430 = ~n1424 & n1429;
  assign n1431 = n1396 & n1430;
  assign n1432 = ~n1395 & ~n1431;
  assign n1433 = n1291 & ~n1432;
  assign n1434 = n1288 ^ n1243;
  assign n1435 = x97 & x108;
  assign n1436 = n1290 & ~n1435;
  assign n1437 = n1436 ^ n1243;
  assign n1438 = n1434 & ~n1437;
  assign n1439 = n1438 ^ n1288;
  assign n1440 = n1233 & n1439;
  assign n1441 = ~n1433 & ~n1440;
  assign n1442 = n1300 & ~n1441;
  assign n1443 = x86 & x94;
  assign n1444 = n1442 & ~n1443;
  assign n1445 = n1444 ^ n1327;
  assign n1446 = ~n1329 & n1445;
  assign n1447 = n1446 ^ n1327;
  assign n1448 = n1304 & ~n1447;
  assign n1449 = n1326 & ~n1448;
  assign n1450 = ~x90 & n1247;
  assign n1451 = x93 ^ x35;
  assign n1452 = n1450 & n1451;
  assign n1453 = ~n1449 & ~n1452;
  assign n1454 = n1286 & ~n1453;
  assign n1455 = ~n1282 & ~n1454;
  assign n1461 = n1460 ^ n1455;
  assign n1462 = n1254 & ~n1461;
  assign n1463 = n1462 ^ n1455;
  assign n1464 = ~n1286 & n1463;
  assign n1465 = x97 & n1306;
  assign n1466 = n1442 & n1465;
  assign n1467 = n1286 & n1306;
  assign n1468 = ~x35 & n1467;
  assign n1469 = n1466 & n1468;
  assign n1470 = ~n1283 & ~n1469;
  assign n1471 = x1091 & x1093;
  assign n1472 = ~x833 & x957;
  assign n1473 = n1471 & n1472;
  assign n1474 = ~x1091 & x1093;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = x950 & x1092;
  assign n1477 = x829 & n1476;
  assign n1478 = n1475 & n1477;
  assign n1479 = ~x841 & n1478;
  assign n1480 = n1247 & n1479;
  assign n1481 = x1093 & n1478;
  assign n1482 = ~x46 & ~x94;
  assign n1483 = x97 ^ x36;
  assign n1484 = n1482 & n1483;
  assign n1485 = n1481 & n1484;
  assign n1486 = ~n1480 & ~n1485;
  assign n1487 = ~n1470 & ~n1486;
  assign n1488 = ~x174 & ~x189;
  assign n1489 = ~x144 & n1488;
  assign n1490 = ~x142 & ~x299;
  assign n1491 = ~n1489 & n1490;
  assign n1492 = ~x152 & ~x166;
  assign n1493 = ~x161 & n1492;
  assign n1494 = ~x146 & x299;
  assign n1495 = ~n1493 & n1494;
  assign n1496 = ~n1491 & ~n1495;
  assign n1497 = ~n1259 & n1496;
  assign n1498 = n1487 & n1497;
  assign n1499 = ~x35 & n1241;
  assign n1500 = ~x97 & ~n1499;
  assign n1501 = ~x137 & ~n1500;
  assign n1502 = ~n1498 & n1501;
  assign n1503 = n1301 & n1303;
  assign n1504 = ~x109 & ~x110;
  assign n1505 = ~n1235 & ~n1504;
  assign n1506 = n1292 & ~n1505;
  assign n1507 = ~n1503 & n1506;
  assign n1508 = n1302 & ~n1507;
  assign n1509 = n1326 & ~n1508;
  assign n1510 = x225 ^ x35;
  assign n1511 = n1510 ^ x225;
  assign n1512 = ~x40 & ~x51;
  assign n1513 = n1248 & n1512;
  assign n1514 = n1513 ^ x225;
  assign n1515 = ~n1511 & n1514;
  assign n1516 = n1515 ^ x225;
  assign n1517 = ~x93 & n1516;
  assign n1518 = n1517 ^ x35;
  assign n1519 = n1450 & ~n1518;
  assign n1520 = ~x95 & ~n1519;
  assign n1521 = ~n1509 & n1520;
  assign n1522 = ~n1449 & n1521;
  assign n1523 = ~n1502 & ~n1522;
  assign n1524 = ~n1464 & n1523;
  assign n1525 = n1524 ^ x234;
  assign n1526 = n1285 & n1525;
  assign n1527 = n1526 ^ x234;
  assign n1528 = ~n1262 & ~n1527;
  assign n1529 = ~x228 & ~n1463;
  assign n1530 = x105 & x228;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~x216 & ~x221;
  assign n1533 = ~x215 & x299;
  assign n1534 = n1532 & n1533;
  assign n1535 = ~n1531 & n1534;
  assign n1536 = ~x223 & ~x224;
  assign n1537 = ~x222 & n1536;
  assign n1538 = ~x299 & n1537;
  assign n1539 = ~n1535 & ~n1538;
  assign n1540 = n1528 & ~n1539;
  assign n1541 = ~x215 & n1532;
  assign n1542 = ~n1531 & n1541;
  assign n1543 = ~x216 & x833;
  assign n1544 = ~x929 & n1543;
  assign n1545 = ~x221 & x265;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~x215 & ~n1546;
  assign n1548 = x221 & ~n1543;
  assign n1549 = ~x215 & ~n1548;
  assign n1550 = ~x1144 & ~n1549;
  assign n1551 = ~n1547 & ~n1550;
  assign n1552 = ~x332 & ~n1551;
  assign n1553 = ~n1541 & ~n1552;
  assign n1554 = x299 & ~n1553;
  assign n1555 = x153 & ~n1530;
  assign n1556 = ~x332 & n1555;
  assign n1557 = n1541 & ~n1556;
  assign n1558 = n1554 & ~n1557;
  assign n1559 = ~n1542 & n1558;
  assign n1560 = ~n1540 & ~n1559;
  assign n1561 = ~x75 & ~x100;
  assign n1562 = ~x74 & n1561;
  assign n1563 = ~x38 & ~x54;
  assign n1564 = n1562 & n1563;
  assign n1565 = ~x87 & ~x92;
  assign n1566 = ~x39 & n1565;
  assign n1567 = n1564 & n1566;
  assign n1568 = ~x56 & ~x62;
  assign n1569 = ~x55 & n1568;
  assign n1570 = ~x57 & ~x59;
  assign n1571 = n1569 & n1570;
  assign n1572 = n1567 & n1571;
  assign n1573 = ~n1560 & n1572;
  assign n1574 = n1254 & n1265;
  assign n1575 = n1567 & n1574;
  assign n1576 = n1570 & n1575;
  assign n1577 = x57 & ~x59;
  assign n1578 = n1568 & n1577;
  assign n1579 = n1575 & n1578;
  assign n1580 = ~x55 & n1579;
  assign n1581 = n1571 & n1574;
  assign n1582 = ~x74 & ~x92;
  assign n1583 = ~x54 & n1582;
  assign n1584 = ~x87 & n1561;
  assign n1585 = n1583 & n1584;
  assign n1586 = x38 & ~x39;
  assign n1587 = n1585 & n1586;
  assign n1588 = n1581 & n1587;
  assign n1589 = ~x39 & ~x87;
  assign n1590 = ~x38 & n1589;
  assign n1591 = ~x92 & n1561;
  assign n1592 = n1590 & n1591;
  assign n1593 = ~x74 & n1592;
  assign n1594 = ~x57 & n1568;
  assign n1595 = x54 & x59;
  assign n1596 = n1594 & ~n1595;
  assign n1597 = ~x54 & ~x59;
  assign n1598 = n1597 ^ x55;
  assign n1599 = n1596 & ~n1598;
  assign n1600 = n1593 & n1599;
  assign n1601 = n1574 & n1600;
  assign n1602 = ~n1588 & ~n1601;
  assign n1603 = ~n1580 & n1602;
  assign n1604 = n1581 & n1590;
  assign n1605 = x74 ^ x54;
  assign n1606 = n1605 ^ x75;
  assign n1607 = n1606 ^ x92;
  assign n1608 = x92 ^ x74;
  assign n1609 = x75 ^ x74;
  assign n1610 = n1608 & n1609;
  assign n1611 = n1610 ^ x74;
  assign n1612 = n1607 & ~n1611;
  assign n1613 = n1604 & n1612;
  assign n1614 = ~x100 & n1613;
  assign n1615 = n1603 & ~n1614;
  assign n1616 = x62 ^ x56;
  assign n1617 = ~x55 & n1616;
  assign n1618 = n1576 & n1617;
  assign n1619 = ~x74 & ~x75;
  assign n1620 = n1563 & n1619;
  assign n1621 = x87 ^ x39;
  assign n1622 = n1621 ^ x92;
  assign n1623 = n1622 ^ x100;
  assign n1624 = x92 ^ x87;
  assign n1625 = x100 ^ x87;
  assign n1626 = n1624 & n1625;
  assign n1627 = n1626 ^ x87;
  assign n1628 = n1623 & ~n1627;
  assign n1629 = n1620 & n1628;
  assign n1630 = n1581 & n1629;
  assign n1631 = ~n1618 & ~n1630;
  assign n1632 = n1615 & n1631;
  assign n1633 = n1576 & ~n1632;
  assign n1634 = ~x228 & n1633;
  assign n1635 = n1541 & n1634;
  assign n1636 = n1541 & ~n1555;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = x234 & n1284;
  assign n1639 = n1530 & ~n1638;
  assign n1640 = ~n1633 & n1639;
  assign n1641 = ~n1618 & ~n1640;
  assign n1642 = ~n1637 & n1641;
  assign n1643 = ~x105 & x228;
  assign n1644 = ~x137 & ~n1643;
  assign n1645 = n1541 & ~n1644;
  assign n1646 = ~x228 & n1570;
  assign n1647 = n1555 & ~n1646;
  assign n1648 = n1645 & ~n1647;
  assign n1649 = ~n1632 & n1648;
  assign n1650 = ~n1553 & ~n1571;
  assign n1651 = ~n1649 & n1650;
  assign n1652 = ~n1642 & n1651;
  assign n1653 = n1564 & n1624;
  assign n1654 = ~n1558 & n1585;
  assign n1655 = ~n1653 & ~n1654;
  assign n1656 = ~x39 & ~n1655;
  assign n1657 = n1563 & n1582;
  assign n1658 = n1584 & n1657;
  assign n1659 = ~n1656 & ~n1658;
  assign n1660 = ~x137 & ~x332;
  assign n1661 = n1538 & n1660;
  assign n1662 = x153 & n1643;
  assign n1663 = n1645 & ~n1662;
  assign n1664 = ~x332 & ~n1663;
  assign n1665 = n1554 & n1664;
  assign n1666 = ~n1661 & ~n1665;
  assign n1667 = ~n1659 & n1666;
  assign n1668 = n1574 & n1667;
  assign n1669 = ~n1567 & n1571;
  assign n1670 = ~n1668 & n1669;
  assign n1671 = ~x146 & ~n1493;
  assign n1672 = ~x210 & ~n1671;
  assign n1673 = n1660 & ~n1672;
  assign n1674 = n1554 & n1673;
  assign n1675 = ~x142 & ~n1489;
  assign n1676 = ~x198 & ~n1675;
  assign n1677 = n1661 & ~n1676;
  assign n1678 = x100 ^ x75;
  assign n1679 = n1583 & n1678;
  assign n1680 = ~n1677 & n1679;
  assign n1681 = x137 & n1561;
  assign n1682 = n1612 & n1681;
  assign n1683 = ~n1680 & ~n1682;
  assign n1684 = ~n1674 & ~n1683;
  assign n1685 = n1574 & n1684;
  assign n1686 = n1590 & n1685;
  assign n1687 = n1686 ^ n1558;
  assign n1688 = n1530 & n1534;
  assign n1689 = ~n1538 & ~n1688;
  assign n1690 = ~x332 & ~n1638;
  assign n1691 = ~n1689 & n1690;
  assign n1692 = n1691 ^ n1686;
  assign n1693 = ~x39 & x252;
  assign n1694 = ~n1653 & n1693;
  assign n1695 = ~n1671 & n1694;
  assign n1696 = ~x228 & n1629;
  assign n1697 = ~n1695 & n1696;
  assign n1698 = n1574 & n1697;
  assign n1699 = n1541 & n1698;
  assign n1700 = n1699 ^ n1686;
  assign n1701 = ~n1686 & n1700;
  assign n1702 = n1701 ^ n1686;
  assign n1703 = ~n1692 & ~n1702;
  assign n1704 = n1703 ^ n1701;
  assign n1705 = n1704 ^ n1686;
  assign n1706 = n1705 ^ n1699;
  assign n1707 = ~n1687 & n1706;
  assign n1708 = n1707 ^ n1686;
  assign n1709 = n1670 & ~n1708;
  assign n1710 = ~x224 & x833;
  assign n1711 = x222 & ~n1710;
  assign n1712 = ~x223 & ~n1711;
  assign n1713 = x1144 & ~n1712;
  assign n1714 = x224 ^ x222;
  assign n1715 = x265 ^ x224;
  assign n1716 = n1715 ^ x265;
  assign n1717 = n1716 ^ n1714;
  assign n1718 = x929 ^ x833;
  assign n1719 = x833 & n1718;
  assign n1720 = n1719 ^ x265;
  assign n1721 = n1720 ^ x833;
  assign n1722 = ~n1717 & n1721;
  assign n1723 = n1722 ^ n1719;
  assign n1724 = n1723 ^ x833;
  assign n1725 = n1714 & n1724;
  assign n1726 = n1725 ^ x222;
  assign n1727 = ~x223 & ~n1726;
  assign n1728 = ~n1713 & ~n1727;
  assign n1729 = ~x299 & n1571;
  assign n1730 = n1728 & n1729;
  assign n1731 = ~n1709 & ~n1730;
  assign n1732 = ~n1652 & n1731;
  assign n1733 = ~n1573 & n1732;
  assign n1734 = ~x332 & ~n1733;
  assign n1735 = ~n1530 & n1541;
  assign n1736 = ~x154 & n1735;
  assign n1737 = ~x215 & x221;
  assign n1738 = n1543 & n1737;
  assign n1739 = x939 & n1738;
  assign n1740 = x216 & ~x221;
  assign n1741 = ~x215 & n1740;
  assign n1742 = x276 & n1741;
  assign n1743 = ~n1739 & ~n1742;
  assign n1744 = ~n1736 & n1743;
  assign n1745 = x1146 & ~n1549;
  assign n1746 = n1744 & ~n1745;
  assign n1747 = n1530 & n1541;
  assign n1748 = n1284 & n1747;
  assign n1749 = x239 & n1748;
  assign n1750 = n1746 & ~n1749;
  assign n1751 = n1541 & ~n1729;
  assign n1752 = ~n1463 & n1572;
  assign n1753 = ~n1633 & ~n1752;
  assign n1754 = ~x228 & ~n1753;
  assign n1755 = n1754 ^ n1729;
  assign n1756 = n1571 & n1698;
  assign n1757 = n1756 ^ n1751;
  assign n1758 = n1755 & n1757;
  assign n1759 = n1758 ^ n1756;
  assign n1760 = n1751 & n1759;
  assign n1761 = n1760 ^ n1729;
  assign n1762 = ~n1750 & ~n1761;
  assign n1763 = n1541 & n1567;
  assign n1764 = x299 & n1763;
  assign n1765 = ~n1285 & n1764;
  assign n1766 = n1529 & n1765;
  assign n1767 = ~n1284 & ~n1567;
  assign n1768 = ~n1285 & ~n1767;
  assign n1769 = ~n1689 & n1768;
  assign n1770 = ~n1766 & ~n1769;
  assign n1771 = x239 & ~n1770;
  assign n1772 = ~x299 & ~n1712;
  assign n1773 = x1146 & n1772;
  assign n1774 = ~x223 & ~x299;
  assign n1775 = x222 & n1774;
  assign n1776 = n1710 & n1775;
  assign n1777 = x939 & n1776;
  assign n1778 = x224 & n1774;
  assign n1779 = ~x222 & n1778;
  assign n1780 = x276 & n1779;
  assign n1781 = ~n1777 & ~n1780;
  assign n1782 = ~n1773 & n1781;
  assign n1783 = ~n1771 & n1782;
  assign n1784 = n1571 & ~n1783;
  assign n1785 = ~n1762 & ~n1784;
  assign n1786 = x274 & n1741;
  assign n1787 = ~x151 & n1735;
  assign n1788 = n1787 ^ n1541;
  assign n1789 = ~n1786 & ~n1788;
  assign n1790 = ~x927 & n1738;
  assign n1791 = n1789 & ~n1790;
  assign n1792 = ~x1145 & ~n1549;
  assign n1793 = n1791 & ~n1792;
  assign n1794 = x235 & n1748;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1761 & ~n1795;
  assign n1797 = x235 & ~n1770;
  assign n1798 = x1145 & n1772;
  assign n1799 = ~x274 & n1779;
  assign n1800 = x927 & n1776;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = ~n1798 & n1801;
  assign n1803 = ~n1797 & n1802;
  assign n1804 = n1571 & ~n1803;
  assign n1805 = ~n1796 & ~n1804;
  assign n1806 = x284 & n1285;
  assign n1807 = n1806 ^ x146;
  assign n1808 = ~n1531 & ~n1807;
  assign n1809 = n1808 ^ x146;
  assign n1810 = n1763 & n1809;
  assign n1811 = ~n1284 & n1747;
  assign n1812 = ~x284 & n1811;
  assign n1813 = ~x264 & n1741;
  assign n1814 = x944 & n1738;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1812 & n1815;
  assign n1817 = x146 & n1735;
  assign n1818 = x1143 & ~n1549;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = n1816 & n1819;
  assign n1821 = ~n1699 & ~n1820;
  assign n1822 = x299 & ~n1821;
  assign n1823 = ~n1530 & ~n1698;
  assign n1824 = x284 & ~n1284;
  assign n1825 = n1541 & ~n1824;
  assign n1826 = ~n1643 & n1825;
  assign n1827 = ~n1823 & n1826;
  assign n1828 = n1822 & ~n1827;
  assign n1829 = ~n1764 & ~n1828;
  assign n1830 = ~n1810 & ~n1829;
  assign n1831 = ~x238 & ~n1770;
  assign n1832 = x284 & n1538;
  assign n1833 = ~n1768 & n1832;
  assign n1834 = x264 & n1779;
  assign n1835 = n1571 & ~n1834;
  assign n1836 = ~x944 & n1776;
  assign n1837 = n1835 & ~n1836;
  assign n1838 = ~x1143 & n1772;
  assign n1839 = n1837 & ~n1838;
  assign n1840 = ~n1833 & n1839;
  assign n1841 = ~n1831 & n1840;
  assign n1842 = ~n1830 & n1841;
  assign n1843 = n1826 ^ n1820;
  assign n1844 = x228 & x238;
  assign n1845 = n1826 & n1844;
  assign n1846 = n1845 ^ n1635;
  assign n1847 = ~n1843 & ~n1846;
  assign n1848 = n1847 ^ n1826;
  assign n1849 = ~n1571 & n1848;
  assign n1850 = ~n1842 & ~n1849;
  assign n1851 = ~x249 & ~n1285;
  assign n1852 = n1538 & n1851;
  assign n1853 = n1543 ^ x932;
  assign n1854 = n1853 ^ x932;
  assign n1855 = x1142 ^ x932;
  assign n1856 = ~n1854 & n1855;
  assign n1857 = n1856 ^ x932;
  assign n1858 = n1857 ^ x216;
  assign n1859 = n1858 ^ n1857;
  assign n1860 = n1857 ^ x277;
  assign n1861 = n1860 ^ n1857;
  assign n1862 = n1859 & ~n1861;
  assign n1863 = n1862 ^ n1857;
  assign n1864 = ~x221 & n1863;
  assign n1865 = n1864 ^ n1857;
  assign n1866 = n1533 & ~n1865;
  assign n1867 = ~n1852 & ~n1866;
  assign n1868 = n1572 & ~n1867;
  assign n1904 = n1531 ^ x172;
  assign n1905 = n1904 ^ x172;
  assign n1906 = x262 ^ x249;
  assign n1907 = n1285 & ~n1906;
  assign n1908 = n1907 ^ x249;
  assign n1909 = n1908 ^ x172;
  assign n1910 = ~n1905 & ~n1909;
  assign n1911 = n1910 ^ x172;
  assign n1869 = ~n1530 & ~n1634;
  assign n1870 = ~n1756 & n1869;
  assign n1871 = ~x262 & ~n1870;
  assign n1872 = n1634 ^ n1284;
  assign n1873 = n1872 ^ n1284;
  assign n1874 = n1284 ^ x172;
  assign n1875 = n1874 ^ n1284;
  assign n1876 = ~n1873 & ~n1875;
  assign n1877 = n1876 ^ n1284;
  assign n1878 = ~n1530 & n1877;
  assign n1879 = n1878 ^ n1284;
  assign n1880 = ~n1871 & ~n1879;
  assign n1881 = n1541 & ~n1880;
  assign n1882 = n1865 ^ x1142;
  assign n1883 = ~x215 & n1882;
  assign n1884 = n1883 ^ x1142;
  assign n1885 = ~n1881 & ~n1884;
  assign n1886 = x262 & n1571;
  assign n1887 = n1699 & n1886;
  assign n1888 = ~x249 & n1284;
  assign n1889 = n1747 & n1888;
  assign n1890 = ~n1729 & ~n1889;
  assign n1891 = ~n1887 & n1890;
  assign n1892 = ~n1885 & n1891;
  assign n1893 = x262 & ~n1768;
  assign n1894 = n1538 & ~n1888;
  assign n1895 = ~n1893 & n1894;
  assign n1896 = x1142 & n1772;
  assign n1897 = ~x277 & n1779;
  assign n1898 = x932 & n1776;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = ~n1896 & n1899;
  assign n1901 = ~n1895 & n1900;
  assign n1902 = n1571 & ~n1901;
  assign n1903 = ~n1892 & ~n1902;
  assign n1912 = n1911 ^ n1903;
  assign n1913 = n1912 ^ n1903;
  assign n1914 = n1903 ^ n1534;
  assign n1915 = n1914 ^ n1903;
  assign n1916 = ~n1913 & n1915;
  assign n1917 = n1916 ^ n1903;
  assign n1918 = n1868 & ~n1917;
  assign n1919 = n1918 ^ n1903;
  assign n1920 = ~x935 & n1738;
  assign n1921 = x270 & n1741;
  assign n1922 = ~n1920 & ~n1921;
  assign n1923 = ~x1141 & ~n1549;
  assign n1924 = n1922 & ~n1923;
  assign n1925 = n1530 ^ x171;
  assign n1926 = n1925 ^ x171;
  assign n1927 = x861 & ~n1284;
  assign n1928 = n1927 ^ x171;
  assign n1929 = n1926 & ~n1928;
  assign n1930 = n1929 ^ x171;
  assign n1931 = n1541 & n1930;
  assign n1932 = n1924 & ~n1931;
  assign n1933 = ~n1542 & ~n1932;
  assign n1934 = n1567 & ~n1933;
  assign n1935 = x299 & ~n1934;
  assign n1936 = ~n1283 & n1927;
  assign n1937 = ~n1539 & ~n1936;
  assign n1938 = ~n1935 & ~n1937;
  assign n1939 = n1927 ^ x299;
  assign n1940 = n1939 ^ n1927;
  assign n1941 = n1932 ^ x861;
  assign n1942 = ~n1699 & n1941;
  assign n1943 = n1942 ^ x861;
  assign n1944 = n1943 ^ n1927;
  assign n1945 = n1940 & n1944;
  assign n1946 = n1945 ^ n1927;
  assign n1947 = ~n1567 & n1946;
  assign n1948 = ~n1938 & ~n1947;
  assign n1949 = ~x1141 & n1772;
  assign n1950 = ~x935 & n1776;
  assign n1951 = x270 & n1779;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1949 & n1952;
  assign n1954 = ~n1948 & n1953;
  assign n1955 = x241 & ~n1770;
  assign n1956 = n1571 & ~n1955;
  assign n1957 = ~n1954 & n1956;
  assign n1958 = ~n1571 & ~n1748;
  assign n1959 = ~x241 & ~n1571;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = n1932 ^ n1635;
  assign n1962 = n1961 ^ n1932;
  assign n1963 = n1941 & n1962;
  assign n1964 = n1963 ^ n1932;
  assign n1965 = ~n1960 & ~n1964;
  assign n1966 = ~n1957 & ~n1965;
  assign n1967 = x1140 & ~n1549;
  assign n1968 = x221 ^ x216;
  assign n1969 = x282 ^ x221;
  assign n1970 = n1969 ^ x282;
  assign n1971 = n1970 ^ n1968;
  assign n1972 = x921 ^ x833;
  assign n1973 = x833 & n1972;
  assign n1974 = n1973 ^ x282;
  assign n1975 = n1974 ^ x833;
  assign n1976 = n1971 & n1975;
  assign n1977 = n1976 ^ n1973;
  assign n1978 = n1977 ^ x833;
  assign n1979 = n1968 & n1978;
  assign n1980 = n1979 ^ x221;
  assign n1981 = ~x215 & ~n1980;
  assign n1982 = ~n1967 & ~n1981;
  assign n1983 = ~x170 & n1735;
  assign n1984 = n1983 ^ n1541;
  assign n1985 = ~n1982 & ~n1984;
  assign n1986 = n1985 ^ x869;
  assign n1987 = n1985 ^ n1811;
  assign n1988 = n1985 ^ n1635;
  assign n1989 = ~n1985 & n1988;
  assign n1990 = n1989 ^ n1985;
  assign n1991 = ~n1987 & ~n1990;
  assign n1992 = n1991 ^ n1989;
  assign n1993 = n1992 ^ n1985;
  assign n1994 = n1993 ^ n1635;
  assign n1995 = n1986 & n1994;
  assign n1996 = n1995 ^ x869;
  assign n1997 = ~n1571 & n1996;
  assign n1999 = x248 & ~n1958;
  assign n1998 = n1571 & n1770;
  assign n2000 = n1999 ^ n1998;
  assign n2001 = n2000 ^ n1999;
  assign n2002 = x299 & ~n1982;
  assign n2003 = n1529 & n1567;
  assign n2004 = n1823 & ~n2003;
  assign n2005 = n2004 ^ x869;
  assign n2006 = n2005 ^ x869;
  assign n2007 = x869 ^ x170;
  assign n2008 = n2006 & ~n2007;
  assign n2009 = n2008 ^ x869;
  assign n2010 = n1541 & ~n2009;
  assign n2011 = n2002 & ~n2010;
  assign n2012 = x1140 & n1772;
  assign n2013 = x869 & ~n1284;
  assign n2014 = n1538 & n2013;
  assign n2015 = ~n2012 & ~n2014;
  assign n2016 = x921 & n1776;
  assign n2017 = ~x282 & n1779;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = n2015 & n2018;
  assign n2020 = ~n2011 & n2019;
  assign n2021 = n2020 ^ n1999;
  assign n2022 = n2001 & ~n2021;
  assign n2023 = n2022 ^ n1999;
  assign n2024 = ~n1997 & ~n2023;
  assign n2025 = x862 ^ x247;
  assign n2026 = ~n1768 & n2025;
  assign n2027 = n2026 ^ x247;
  assign n2028 = n1538 & ~n2027;
  assign n2029 = x148 & n1735;
  assign n2030 = ~x920 & n1738;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~x1139 & ~n1549;
  assign n2033 = x281 & n1741;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = n2031 & n2034;
  assign n2036 = n1284 ^ x862;
  assign n2037 = n2036 ^ x862;
  assign n2038 = n2025 & n2037;
  assign n2039 = n2038 ^ x862;
  assign n2040 = n1747 & ~n2039;
  assign n2041 = n2035 & ~n2040;
  assign n2042 = ~n1763 & ~n2041;
  assign n2043 = n2042 ^ x862;
  assign n2044 = ~n1699 & ~n2043;
  assign n2045 = n2044 ^ x862;
  assign n2046 = x299 & ~n2045;
  assign n2047 = x281 & n1779;
  assign n2048 = n1571 & ~n2047;
  assign n2049 = ~x920 & n1776;
  assign n2050 = n2048 & ~n2049;
  assign n2051 = ~x1139 & n1772;
  assign n2052 = n2050 & ~n2051;
  assign n2053 = ~n2046 & n2052;
  assign n2054 = ~n2028 & n2053;
  assign n2055 = n1531 ^ x148;
  assign n2056 = n2055 ^ x148;
  assign n2057 = n1285 & n2025;
  assign n2058 = n2057 ^ x247;
  assign n2059 = n2058 ^ x148;
  assign n2060 = ~n2056 & ~n2059;
  assign n2061 = n2060 ^ x148;
  assign n2062 = n1764 & n2061;
  assign n2063 = n2054 & ~n2062;
  assign n2064 = n2041 ^ x862;
  assign n2065 = n1635 ^ x862;
  assign n2066 = n2065 ^ x862;
  assign n2067 = n2064 & ~n2066;
  assign n2068 = n2067 ^ x862;
  assign n2069 = ~n1571 & n2068;
  assign n2070 = ~n2063 & ~n2069;
  assign n2071 = ~x1138 & ~n1549;
  assign n2072 = x269 & n1741;
  assign n2073 = ~x940 & n1738;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = ~n2071 & n2074;
  assign n2076 = x299 & n2075;
  assign n2077 = x877 ^ x246;
  assign n2078 = n1285 & n2077;
  assign n2079 = n2078 ^ x246;
  assign n2080 = n2079 ^ x169;
  assign n2081 = ~n1531 & ~n2080;
  assign n2082 = n2081 ^ x169;
  assign n2083 = n2082 ^ n1567;
  assign n2084 = n2083 ^ n2082;
  assign n2085 = x877 & ~n1284;
  assign n2086 = n2085 ^ x169;
  assign n2087 = ~n1823 & ~n2086;
  assign n2088 = n2087 ^ x169;
  assign n2089 = n2088 ^ n2082;
  assign n2090 = ~n2084 & n2089;
  assign n2091 = n2090 ^ n2082;
  assign n2092 = n1541 & n2091;
  assign n2093 = n2076 & ~n2092;
  assign n2094 = x1138 & n1772;
  assign n2095 = ~x269 & n1779;
  assign n2096 = x877 & n1538;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = ~n2094 & n2097;
  assign n2099 = x940 & n1776;
  assign n2100 = n2098 & ~n2099;
  assign n2101 = n2100 ^ x246;
  assign n2102 = ~n1769 & ~n2101;
  assign n2103 = n2102 ^ x246;
  assign n2104 = n1571 & ~n2103;
  assign n2105 = ~n2093 & n2104;
  assign n2106 = n1869 ^ x169;
  assign n2107 = n2106 ^ x169;
  assign n2108 = ~n2086 & ~n2107;
  assign n2109 = n2108 ^ x169;
  assign n2110 = n1541 & n2109;
  assign n2111 = n2075 & ~n2110;
  assign n2112 = x246 & n1748;
  assign n2113 = ~n1571 & ~n2112;
  assign n2114 = ~n2111 & n2113;
  assign n2115 = ~n2105 & ~n2114;
  assign n2158 = n1635 ^ x878;
  assign n2159 = n2158 ^ x878;
  assign n2121 = ~x280 & n1741;
  assign n2122 = n1530 ^ x168;
  assign n2123 = n2122 ^ x168;
  assign n2124 = x878 & ~n1284;
  assign n2125 = n2124 ^ x168;
  assign n2126 = n2123 & ~n2125;
  assign n2127 = n2126 ^ x168;
  assign n2128 = n1541 & ~n2127;
  assign n2129 = ~n2121 & ~n2128;
  assign n2117 = x1137 & ~n1549;
  assign n2118 = x933 & n1738;
  assign n2119 = ~n2117 & ~n2118;
  assign n2160 = x240 & n1748;
  assign n2161 = n2119 & ~n2160;
  assign n2162 = n2129 & n2161;
  assign n2163 = n2162 ^ x878;
  assign n2164 = ~n2159 & ~n2163;
  assign n2165 = n2164 ^ x878;
  assign n2116 = n1567 & n1769;
  assign n2120 = x299 & n2119;
  assign n2130 = n2129 ^ n1699;
  assign n2131 = n2130 ^ n2129;
  assign n2132 = n2129 ^ x878;
  assign n2133 = n2131 & ~n2132;
  assign n2134 = n2133 ^ n2129;
  assign n2135 = n2120 & n2134;
  assign n2136 = ~n2116 & ~n2135;
  assign n2137 = ~n1764 & n2136;
  assign n2138 = ~n1567 & ~n1769;
  assign n2139 = n1534 & ~n2138;
  assign n2140 = x878 ^ x240;
  assign n2141 = n1285 & n2140;
  assign n2142 = n2141 ^ x240;
  assign n2143 = n2142 ^ n1531;
  assign n2144 = n2143 ^ n2142;
  assign n2145 = n2142 ^ x168;
  assign n2146 = n2144 & ~n2145;
  assign n2147 = n2146 ^ n2142;
  assign n2148 = n2139 & n2147;
  assign n2149 = ~n2137 & ~n2148;
  assign n2150 = ~x1137 & n1772;
  assign n2151 = n1538 & ~n2124;
  assign n2152 = x280 & n1779;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2150 & n2153;
  assign n2155 = ~x933 & n1776;
  assign n2156 = n2154 & ~n2155;
  assign n2157 = ~n2149 & n2156;
  assign n2166 = n2165 ^ n2157;
  assign n2167 = n2166 ^ n2165;
  assign n2168 = x240 & n1538;
  assign n2169 = n1768 & n2168;
  assign n2170 = n2169 ^ n2165;
  assign n2171 = n2170 ^ n2165;
  assign n2172 = ~n2167 & ~n2171;
  assign n2173 = n2172 ^ n2165;
  assign n2174 = n1571 & ~n2173;
  assign n2175 = n2174 ^ n2165;
  assign n2176 = n1531 & n1571;
  assign n2177 = x875 & ~n1284;
  assign n2178 = n2177 ^ x166;
  assign n2179 = ~n1823 & n2178;
  assign n2180 = n2179 ^ x166;
  assign n2181 = n2176 & ~n2180;
  assign n2182 = n1541 & ~n2181;
  assign n2183 = ~x875 & ~n1284;
  assign n2184 = n2183 ^ x166;
  assign n2185 = ~n1869 & ~n2184;
  assign n2186 = n2185 ^ x166;
  assign n2187 = ~n1572 & ~n2186;
  assign n2188 = n2187 ^ n1531;
  assign n2189 = n2187 ^ n1571;
  assign n2190 = n2189 ^ n1571;
  assign n2191 = ~n1572 & n2180;
  assign n2192 = x875 ^ x245;
  assign n2193 = n1285 & n2192;
  assign n2194 = n2193 ^ x245;
  assign n2195 = ~n2191 & ~n2194;
  assign n2196 = n2195 ^ n1571;
  assign n2197 = ~n2190 & n2196;
  assign n2198 = n2197 ^ n1571;
  assign n2199 = ~n2188 & ~n2198;
  assign n2200 = n2199 ^ n1531;
  assign n2201 = n2182 & n2200;
  assign n2202 = x1136 & ~n1549;
  assign n2203 = x928 & n1738;
  assign n2204 = x266 & n1741;
  assign n2205 = ~n2203 & ~n2204;
  assign n2206 = ~n2202 & n2205;
  assign n2207 = ~n1729 & n2206;
  assign n2208 = ~n2201 & n2207;
  assign n2209 = ~x1136 & n1772;
  assign n2210 = ~x266 & n1779;
  assign n2211 = ~x928 & n1776;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2209 & n2212;
  assign n2214 = n1571 & ~n2213;
  assign n2215 = n1538 & n1571;
  assign n2216 = n1768 ^ x875;
  assign n2217 = n2216 ^ x875;
  assign n2218 = n2192 & n2217;
  assign n2219 = n2218 ^ x875;
  assign n2220 = n2215 & ~n2219;
  assign n2221 = ~n2214 & ~n2220;
  assign n2222 = ~n2208 & n2221;
  assign n2223 = x244 & ~n1770;
  assign n2224 = x879 & ~n1768;
  assign n2225 = n1534 & ~n1823;
  assign n2226 = ~n1538 & ~n2225;
  assign n2227 = n2224 & ~n2226;
  assign n2228 = x279 & n1779;
  assign n2229 = n1571 & ~n2228;
  assign n2230 = x938 & n1776;
  assign n2231 = n2229 & ~n2230;
  assign n2232 = x1135 & n1772;
  assign n2233 = n2231 & ~n2232;
  assign n2234 = ~n2227 & n2233;
  assign n2235 = ~n2223 & n2234;
  assign n2236 = n2004 ^ x161;
  assign n2237 = n2236 ^ x161;
  assign n2238 = n2224 ^ x161;
  assign n2239 = ~n2237 & n2238;
  assign n2240 = n2239 ^ x161;
  assign n2241 = n1541 & n2240;
  assign n2242 = n2235 & ~n2241;
  assign n2243 = x879 ^ x244;
  assign n2244 = ~n1284 & n2243;
  assign n2245 = n2244 ^ x244;
  assign n2246 = n2245 ^ x161;
  assign n2247 = ~n1869 & n2246;
  assign n2248 = n2247 ^ x161;
  assign n2249 = n1541 & n2248;
  assign n2250 = ~n1571 & ~n2249;
  assign n2251 = ~n2242 & ~n2250;
  assign n2252 = x1135 & ~n1549;
  assign n2253 = x938 & n1738;
  assign n2254 = x279 & n1741;
  assign n2255 = ~n2253 & ~n2254;
  assign n2256 = ~n2252 & n2255;
  assign n2257 = ~n2251 & n2256;
  assign n2258 = ~x299 & n2235;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = x846 ^ x242;
  assign n2261 = ~n1768 & n2260;
  assign n2262 = n2261 ^ x242;
  assign n2263 = n1538 & ~n2262;
  assign n2264 = ~x930 & n1776;
  assign n2265 = ~x278 & n1779;
  assign n2266 = ~n2264 & ~n2265;
  assign n2267 = n1571 & n2266;
  assign n2268 = ~n2263 & n2267;
  assign n2269 = n2004 ^ x152;
  assign n2270 = n2269 ^ x152;
  assign n2271 = n2262 ^ x152;
  assign n2272 = ~n2270 & n2271;
  assign n2273 = n2272 ^ x152;
  assign n2274 = n1541 & ~n2273;
  assign n2275 = n2268 & ~n2274;
  assign n2276 = n1869 ^ x152;
  assign n2277 = n2276 ^ x152;
  assign n2278 = ~n1284 & n2260;
  assign n2279 = n2278 ^ x242;
  assign n2280 = n2279 ^ x152;
  assign n2281 = ~n2277 & n2280;
  assign n2282 = n2281 ^ x152;
  assign n2283 = n1541 & ~n2282;
  assign n2284 = ~n1571 & ~n2283;
  assign n2285 = ~n2275 & ~n2284;
  assign n2286 = ~x278 & n1741;
  assign n2287 = ~x930 & n1738;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2285 & n2288;
  assign n2290 = ~x299 & n2268;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = n1772 ^ n1549;
  assign n2293 = n1729 & ~n2292;
  assign n2294 = n2293 ^ n1549;
  assign n2295 = ~x1134 & ~n2294;
  assign n2296 = ~n2291 & ~n2295;
  assign n2297 = n1233 & n1244;
  assign n2298 = n1326 & ~n2297;
  assign n2299 = n1444 & n2298;
  assign n2300 = x93 & x841;
  assign n2301 = n1452 & ~n2300;
  assign n2302 = n1513 & ~n2301;
  assign n2303 = ~n1509 & n2302;
  assign n2304 = ~n2299 & n2303;
  assign n2305 = ~n1464 & ~n2304;
  assign n2306 = ~n1255 & ~n2305;
  assign n2307 = n1255 & ~n1260;
  assign n2308 = x32 & ~n2307;
  assign n2309 = ~x70 & ~x95;
  assign n2310 = n1241 & n2309;
  assign n2311 = ~n2308 & n2310;
  assign n2312 = x32 & ~n2311;
  assign n2313 = n1572 & ~n1574;
  assign n2314 = ~n2312 & n2313;
  assign n2315 = ~n2306 & n2314;
  assign n2316 = ~x250 & ~n1496;
  assign n2317 = x824 & n1476;
  assign n2318 = ~x1093 & n2317;
  assign n2319 = ~x1093 & n1477;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = n2316 & ~n2320;
  assign n2322 = ~x41 & ~x101;
  assign n2323 = ~x99 & n2322;
  assign n2324 = ~x113 & n2323;
  assign n2325 = ~x43 & ~x44;
  assign n2326 = ~x42 & ~x114;
  assign n2327 = n2325 & n2326;
  assign n2328 = ~x115 & ~x116;
  assign n2329 = n2327 & n2328;
  assign n2330 = n2324 & n2329;
  assign n2331 = ~x52 & n2330;
  assign n2332 = ~x129 & x250;
  assign n2333 = x683 & ~n2332;
  assign n2334 = ~n2331 & n2333;
  assign n2335 = n2334 ^ n1496;
  assign n2336 = n2335 ^ n2334;
  assign n2337 = n2334 ^ x252;
  assign n2338 = n2336 & n2337;
  assign n2339 = n2338 ^ n2334;
  assign n2340 = ~n2321 & n2339;
  assign n2341 = x100 & ~n2340;
  assign n2342 = ~x87 & x100;
  assign n2343 = ~n1590 & ~n2342;
  assign n2344 = ~x74 & ~n2343;
  assign n2345 = ~n2341 & n2344;
  assign n2380 = ~x979 & ~x984;
  assign n2381 = ~x287 & n2380;
  assign n2382 = ~x252 & ~x1001;
  assign n2383 = x835 & ~n2382;
  assign n2384 = n2381 & n2383;
  assign n2346 = ~x332 & ~x468;
  assign n2354 = ~x969 & ~x971;
  assign n2355 = ~x974 & ~x977;
  assign n2356 = n2354 & n2355;
  assign n2357 = ~x587 & ~x602;
  assign n2358 = ~x961 & ~x967;
  assign n2359 = n2357 & n2358;
  assign n2360 = n2356 & n2359;
  assign n2347 = ~x614 & ~x616;
  assign n2348 = ~x642 & n2347;
  assign n2349 = x603 & n2348;
  assign n2350 = ~x661 & ~x662;
  assign n2351 = ~x681 & n2350;
  assign n2352 = x680 & n2351;
  assign n2353 = ~n2349 & ~n2352;
  assign n2361 = n2360 ^ n2353;
  assign n2362 = n2346 & n2361;
  assign n2363 = n2362 ^ n2353;
  assign n2387 = x299 & n2346;
  assign n2388 = n2363 & ~n2387;
  assign n2389 = ~n1473 & n2317;
  assign n2390 = ~n1478 & ~n2389;
  assign n2391 = ~n2388 & ~n2390;
  assign n2392 = n2384 & n2391;
  assign n2393 = ~n1533 & ~n1774;
  assign n2394 = n2392 & n2393;
  assign n2368 = ~x970 & ~x972;
  assign n2369 = ~x975 & ~x978;
  assign n2370 = n2368 & n2369;
  assign n2371 = ~x907 & ~x947;
  assign n2372 = ~x960 & ~x963;
  assign n2373 = n2371 & n2372;
  assign n2374 = n2370 & n2373;
  assign n2395 = n2346 & n2374;
  assign n2396 = x299 & n2395;
  assign n2397 = n2394 & ~n2396;
  assign n2364 = x224 & n1775;
  assign n2365 = ~n2363 & n2364;
  assign n2366 = x299 & n1737;
  assign n2367 = x216 & n2366;
  assign n2375 = n2374 ^ n2353;
  assign n2376 = n2346 & n2375;
  assign n2377 = n2376 ^ n2353;
  assign n2378 = n2367 & ~n2377;
  assign n2379 = ~n2365 & ~n2378;
  assign n2385 = n1481 & n2384;
  assign n2386 = ~n2379 & n2385;
  assign n2398 = n2397 ^ n2386;
  assign n2399 = n2386 ^ x39;
  assign n2400 = ~n2386 & ~n2399;
  assign n2401 = n2400 ^ n2386;
  assign n2402 = n2398 & ~n2401;
  assign n2403 = n2402 ^ n2400;
  assign n2404 = n2403 ^ n2386;
  assign n2405 = n2404 ^ x39;
  assign n2406 = ~n2345 & ~n2405;
  assign n2407 = n2406 ^ n2345;
  assign n2408 = ~n1632 & ~n2407;
  assign n2409 = ~n1580 & ~n1618;
  assign n2410 = ~n2408 & n2409;
  assign n2411 = ~n2315 & n2410;
  assign n2412 = n1286 & n1572;
  assign n2413 = n1509 & n2412;
  assign n2414 = ~n1752 & ~n2413;
  assign n2415 = n1385 ^ n1214;
  assign n2416 = n1214 ^ x67;
  assign n2417 = n2416 ^ n1214;
  assign n2418 = n2415 & ~n2417;
  assign n2419 = n2418 ^ n1214;
  assign n2420 = n1217 & n2419;
  assign n2421 = n1333 & n2420;
  assign n2422 = ~x85 & n1392;
  assign n2423 = ~n1381 & n2422;
  assign n2424 = ~n2421 & n2423;
  assign n2425 = ~x82 & n2424;
  assign n2426 = ~n2297 & n2425;
  assign n2427 = ~x58 & n1303;
  assign n2428 = ~n2426 & n2427;
  assign n2429 = n2302 & n2428;
  assign n2430 = x103 & ~x314;
  assign n2431 = ~x109 & ~n2430;
  assign n2432 = ~n2429 & n2431;
  assign n2433 = ~n2414 & ~n2432;
  assign n2434 = ~x72 & ~n2433;
  assign n2435 = ~n1455 & n1572;
  assign n2436 = n1256 & n1260;
  assign n2437 = n1225 & n1399;
  assign n2438 = n1246 & n2437;
  assign n2439 = n1220 & n2438;
  assign n2440 = ~x73 & n1253;
  assign n2441 = n2439 & n2440;
  assign n2442 = ~x32 & n1284;
  assign n2443 = n2441 & n2442;
  assign n2444 = n1250 & n1264;
  assign n2445 = ~x58 & x841;
  assign n2446 = n1315 & ~n2445;
  assign n2447 = n2444 & n2446;
  assign n2448 = ~n2443 & ~n2447;
  assign n2449 = ~n2436 & n2448;
  assign n2450 = ~n1265 & n2449;
  assign n2451 = n1250 & n1572;
  assign n2452 = n1326 & n2451;
  assign n2453 = ~n2450 & n2452;
  assign n2454 = ~n2435 & ~n2453;
  assign n2455 = ~n2434 & ~n2454;
  assign n2456 = x158 & x159;
  assign n2457 = x197 & n2456;
  assign n2458 = x160 & x232;
  assign n2459 = n2457 & n2458;
  assign n2460 = x299 & ~n2459;
  assign n2461 = n2346 & ~n2460;
  assign n2462 = x109 & x145;
  assign n2463 = x180 & x181;
  assign n2464 = n2462 & n2463;
  assign n2465 = x182 & x232;
  assign n2466 = n2464 & n2465;
  assign n2467 = x109 & x299;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = n2461 & ~n2468;
  assign n2470 = n2455 & ~n2469;
  assign n2471 = ~x228 & n2470;
  assign n2472 = n1583 & n1604;
  assign n2473 = ~x75 & x100;
  assign n2474 = n2340 & n2473;
  assign n2475 = n2472 & n2474;
  assign n2476 = n1615 & ~n2475;
  assign n2477 = x1093 & n2389;
  assign n2478 = x829 & x1092;
  assign n2479 = ~n1474 & n2478;
  assign n2480 = n2477 & ~n2479;
  assign n2481 = n2384 & n2480;
  assign n2482 = ~n1775 & ~n2366;
  assign n2483 = n2481 & ~n2482;
  assign n2484 = ~n2364 & ~n2367;
  assign n2485 = n2385 & ~n2484;
  assign n2486 = ~n2483 & ~n2485;
  assign n2487 = x39 & n1658;
  assign n2488 = ~n2486 & n2487;
  assign n2489 = n1574 & n2488;
  assign n2490 = ~x228 & ~n2489;
  assign n2491 = n2476 & n2490;
  assign n2492 = ~x30 & x228;
  assign n2493 = n1571 & ~n2492;
  assign n2494 = ~n2491 & n2493;
  assign n2495 = ~n2471 & ~n2494;
  assign n2496 = ~x299 & n2346;
  assign n2497 = ~n2495 & n2496;
  assign n2498 = x602 & n2497;
  assign n2499 = ~x228 & n2455;
  assign n2500 = ~x228 & n1615;
  assign n2501 = ~n1571 & ~n2492;
  assign n2502 = ~n2500 & n2501;
  assign n2503 = ~n2494 & ~n2502;
  assign n2504 = ~n2499 & n2503;
  assign n2505 = ~x299 & ~n2501;
  assign n2506 = x109 & ~x228;
  assign n2507 = n2459 & n2506;
  assign n2508 = n2346 & ~n2507;
  assign n2509 = ~n2505 & n2508;
  assign n2510 = x907 & n2509;
  assign n2511 = ~n2346 & n2352;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = ~n2504 & ~n2512;
  assign n2514 = ~n2498 & ~n2513;
  assign n2515 = ~n2495 & ~n2496;
  assign n2516 = ~n2502 & ~n2515;
  assign n2517 = n2349 ^ x947;
  assign n2518 = ~n2346 & n2517;
  assign n2519 = n2518 ^ x947;
  assign n2520 = ~n2516 & n2519;
  assign n2521 = x587 & n2497;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = x967 & n2497;
  assign n2524 = ~n2504 & n2509;
  assign n2525 = x970 & n2524;
  assign n2526 = ~n2523 & ~n2525;
  assign n2527 = x299 & x972;
  assign n2528 = ~x109 & n2527;
  assign n2529 = ~x299 & x961;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = ~n2466 & ~n2530;
  assign n2532 = ~n2459 & n2527;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n2499 & ~n2533;
  assign n2535 = ~n2527 & ~n2529;
  assign n2536 = n2494 & ~n2535;
  assign n2537 = x972 & n2502;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = ~n2534 & n2538;
  assign n2540 = n2346 & ~n2539;
  assign n2541 = x977 & n2497;
  assign n2542 = x960 & n2524;
  assign n2543 = ~n2541 & ~n2542;
  assign n2544 = x969 & n2497;
  assign n2545 = x963 & n2524;
  assign n2546 = ~n2544 & ~n2545;
  assign n2547 = x971 & n2497;
  assign n2548 = x975 & n2524;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = x974 & n2497;
  assign n2551 = x978 & n2524;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = ~x96 & n1265;
  assign n2554 = ~x90 & ~x93;
  assign n2555 = ~x35 & ~x70;
  assign n2556 = n2554 & n2555;
  assign n2557 = n2553 & n2556;
  assign n2558 = n1246 & n2557;
  assign n2559 = n1229 & n2558;
  assign n2560 = ~x92 & n1564;
  assign n2561 = n1571 & n2560;
  assign n2562 = n2559 & n2561;
  assign n2563 = x39 & ~x72;
  assign n2564 = n2562 & n2563;
  assign n2565 = ~x51 & ~x87;
  assign n2566 = n1232 & n2565;
  assign n2567 = n2564 & n2566;
  assign n2568 = ~n1729 & n1737;
  assign n2569 = ~n2377 & n2568;
  assign n2570 = n1571 & n1775;
  assign n2571 = ~n2363 & n2570;
  assign n2572 = ~n2569 & ~n2571;
  assign n2573 = n2481 & ~n2572;
  assign n2574 = ~n2386 & ~n2573;
  assign n2575 = n2567 & ~n2574;
  assign n2576 = n2476 & ~n2575;
  assign n2577 = ~n2470 & n2576;
  assign n2578 = n2577 ^ x24;
  assign n2579 = ~x954 & n2578;
  assign n2580 = n2579 ^ x24;
  assign n2581 = n1496 & n1694;
  assign n2582 = n1630 & ~n2581;
  assign n2583 = n1753 & ~n2582;
  assign n2584 = n2583 ^ x105;
  assign n2585 = ~x228 & ~n2584;
  assign n2586 = n2585 ^ x105;
  assign n2587 = ~x119 & ~x228;
  assign n2588 = x252 & ~x468;
  assign n2589 = n2587 & n2588;
  assign n2590 = x119 & ~x468;
  assign n2591 = ~x1056 & n2590;
  assign n2592 = ~n2589 & ~n2591;
  assign n2593 = ~x1077 & n2590;
  assign n2594 = ~n2589 & ~n2593;
  assign n2595 = ~x1073 & n2590;
  assign n2596 = ~n2589 & ~n2595;
  assign n2597 = ~x1041 & n2590;
  assign n2598 = ~n2589 & ~n2597;
  assign n2599 = n1249 & n1449;
  assign n2600 = x98 & n2599;
  assign n2601 = x90 ^ x51;
  assign n2602 = n2601 ^ x93;
  assign n2603 = x93 ^ x90;
  assign n2604 = x841 ^ x90;
  assign n2605 = n2603 & n2604;
  assign n2606 = n2605 ^ x90;
  assign n2607 = n2602 & ~n2606;
  assign n2608 = n2555 & n2607;
  assign n2609 = n1247 & n2608;
  assign n2610 = ~n2600 & ~n2609;
  assign n2611 = ~x96 & n2610;
  assign n2612 = ~x98 & x1091;
  assign n2613 = n2320 & ~n2612;
  assign n2614 = ~x72 & ~n2613;
  assign n2615 = ~n2390 & n2614;
  assign n2616 = ~n2611 & n2615;
  assign n2617 = x91 & n1503;
  assign n2618 = ~x24 & ~x58;
  assign n2619 = n2617 & n2618;
  assign n2620 = ~n1466 & ~n2619;
  assign n2621 = ~x122 & n1481;
  assign n2622 = ~x72 & n1249;
  assign n2623 = n1252 & n2622;
  assign n2624 = n2621 & n2623;
  assign n2625 = ~n2620 & n2624;
  assign n2626 = ~n2616 & ~n2625;
  assign n2627 = n1249 & n1263;
  assign n2628 = ~x122 & x829;
  assign n2629 = ~x841 & n2628;
  assign n2630 = n1265 & n2629;
  assign n2631 = n2627 & n2630;
  assign n2632 = ~n2553 & ~n2631;
  assign n2633 = ~n2626 & ~n2632;
  assign n2634 = ~x39 & ~x72;
  assign n2635 = n2553 & n2634;
  assign n2636 = ~n2610 & n2635;
  assign n2637 = ~x87 & ~n2636;
  assign n2638 = ~n2390 & ~n2637;
  assign n2639 = x100 ^ x39;
  assign n2640 = ~x75 & ~n2639;
  assign n2641 = ~n2638 & n2640;
  assign n2642 = ~n2633 & n2641;
  assign n2643 = x232 & n2346;
  assign n2644 = n1489 ^ x299;
  assign n2645 = n2644 ^ n1489;
  assign n2646 = n1493 ^ n1489;
  assign n2647 = n2645 & n2646;
  assign n2648 = n2647 ^ n1489;
  assign n2649 = n2643 & n2648;
  assign n2650 = ~n2331 & ~n2649;
  assign n2651 = x252 & n2650;
  assign n2652 = ~x24 & ~x100;
  assign n2653 = ~x87 & n2652;
  assign n2654 = n2621 & n2653;
  assign n2655 = n2651 & n2654;
  assign n2656 = n1574 & n2655;
  assign n2657 = x75 & ~n2656;
  assign n2658 = ~x39 & ~x100;
  assign n2659 = n1657 & n2658;
  assign n2660 = n1574 & n2659;
  assign n2661 = ~n2657 & n2660;
  assign n2662 = ~n1775 & ~n1778;
  assign n2663 = ~n2363 & ~n2662;
  assign n2664 = ~n1532 & n1533;
  assign n2665 = ~n2377 & n2664;
  assign n2666 = ~n2663 & ~n2665;
  assign n2667 = ~x224 & n1775;
  assign n2668 = ~x216 & n2366;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2666 & ~n2669;
  assign n2671 = n2385 & n2670;
  assign n2672 = x39 & ~n2671;
  assign n2673 = n2621 & n2650;
  assign n2674 = x228 & n2673;
  assign n2675 = x100 & ~n2674;
  assign n2676 = n1565 & n1620;
  assign n2677 = ~n2675 & n2676;
  assign n2678 = ~n2672 & n2677;
  assign n2679 = n1574 & n2678;
  assign n2680 = ~n1567 & ~n2679;
  assign n2681 = ~n2661 & n2680;
  assign n2687 = x335 ^ x334;
  assign n2688 = n2687 ^ x333;
  assign n2685 = x463 ^ x413;
  assign n2683 = x407 ^ x393;
  assign n2682 = x392 ^ x391;
  assign n2684 = n2683 ^ n2682;
  assign n2686 = n2685 ^ n2684;
  assign n2689 = n2688 ^ n2686;
  assign n2690 = x1197 & n2689;
  assign n2696 = x394 ^ x329;
  assign n2697 = n2696 ^ x328;
  assign n2694 = x399 ^ x398;
  assign n2692 = x408 ^ x400;
  assign n2691 = x396 ^ x395;
  assign n2693 = n2692 ^ n2691;
  assign n2695 = n2694 ^ n2693;
  assign n2698 = n2697 ^ n2695;
  assign n2699 = x1198 & n2698;
  assign n2700 = ~n2690 & ~n2699;
  assign n2701 = ~x592 & ~n2700;
  assign n2702 = x591 & ~n2701;
  assign n2703 = ~x590 & ~x592;
  assign n2709 = x390 ^ x324;
  assign n2710 = n2709 ^ x319;
  assign n2707 = x456 ^ x412;
  assign n2705 = x404 ^ x397;
  assign n2704 = x411 ^ x410;
  assign n2706 = n2705 ^ n2704;
  assign n2708 = n2707 ^ n2706;
  assign n2711 = n2710 ^ n2708;
  assign n2712 = x1196 & n2711;
  assign n2718 = x326 ^ x325;
  assign n2719 = n2718 ^ x318;
  assign n2716 = x405 ^ x403;
  assign n2714 = x409 ^ x406;
  assign n2713 = x402 ^ x401;
  assign n2715 = n2714 ^ n2713;
  assign n2717 = n2716 ^ n2715;
  assign n2720 = n2719 ^ n2717;
  assign n2721 = x1199 & n2720;
  assign n2722 = ~n2712 & ~n2721;
  assign n2723 = n2703 & ~n2722;
  assign n2724 = x567 & n2723;
  assign n2725 = n2702 & ~n2724;
  assign n2731 = x371 ^ x370;
  assign n2732 = n2731 ^ x369;
  assign n2729 = x442 ^ x440;
  assign n2727 = x384 ^ x375;
  assign n2726 = x374 ^ x373;
  assign n2728 = n2727 ^ n2726;
  assign n2730 = n2729 ^ n2728;
  assign n2733 = n2732 ^ n2730;
  assign n2734 = x1198 & n2733;
  assign n2740 = x339 ^ x338;
  assign n2741 = n2740 ^ x337;
  assign n2738 = x388 ^ x387;
  assign n2736 = x372 ^ x363;
  assign n2735 = x386 ^ x380;
  assign n2737 = n2736 ^ n2735;
  assign n2739 = n2738 ^ n2737;
  assign n2742 = n2741 ^ n2739;
  assign n2743 = x1196 & n2742;
  assign n2744 = ~n2734 & ~n2743;
  assign n2750 = x365 ^ x364;
  assign n2751 = n2750 ^ x336;
  assign n2748 = x447 ^ x389;
  assign n2746 = x383 ^ x368;
  assign n2745 = x367 ^ x366;
  assign n2747 = n2746 ^ n2745;
  assign n2749 = n2748 ^ n2747;
  assign n2752 = n2751 ^ n2749;
  assign n2753 = x1197 & n2752;
  assign n2754 = n2744 & ~n2753;
  assign n2760 = x377 ^ x376;
  assign n2761 = n2760 ^ x317;
  assign n2758 = x382 ^ x381;
  assign n2756 = x439 ^ x385;
  assign n2755 = x379 ^ x378;
  assign n2757 = n2756 ^ n2755;
  assign n2759 = n2758 ^ n2757;
  assign n2762 = n2761 ^ n2759;
  assign n2763 = x1199 & n2762;
  assign n2764 = ~x591 & ~n2763;
  assign n2765 = n2754 & n2764;
  assign n2766 = ~x590 & ~n2765;
  assign n2772 = x353 ^ x352;
  assign n2773 = n2772 ^ x351;
  assign n2770 = x462 ^ x461;
  assign n2768 = x360 ^ x357;
  assign n2767 = x356 ^ x354;
  assign n2769 = n2768 ^ n2767;
  assign n2771 = n2770 ^ n2769;
  assign n2774 = n2773 ^ n2771;
  assign n2775 = x1199 & n2774;
  assign n2781 = x355 ^ x342;
  assign n2782 = n2781 ^ x320;
  assign n2779 = x455 ^ x452;
  assign n2777 = x460 ^ x458;
  assign n2776 = x441 ^ x361;
  assign n2778 = n2777 ^ n2776;
  assign n2780 = n2779 ^ n2778;
  assign n2783 = n2782 ^ n2780;
  assign n2784 = x1196 & n2783;
  assign n2785 = ~n2775 & ~n2784;
  assign n2791 = x321 ^ x316;
  assign n2792 = n2791 ^ x315;
  assign n2789 = x349 ^ x348;
  assign n2787 = x359 ^ x350;
  assign n2786 = x347 ^ x322;
  assign n2788 = n2787 ^ n2786;
  assign n2790 = n2789 ^ n2788;
  assign n2793 = n2792 ^ n2790;
  assign n2794 = x1198 & n2793;
  assign n2800 = x343 ^ x327;
  assign n2801 = n2800 ^ x323;
  assign n2798 = x450 ^ x362;
  assign n2796 = x358 ^ x346;
  assign n2795 = x345 ^ x344;
  assign n2797 = n2796 ^ n2795;
  assign n2799 = n2798 ^ n2797;
  assign n2802 = n2801 ^ n2799;
  assign n2803 = x1197 & n2802;
  assign n2804 = ~n2794 & ~n2803;
  assign n2805 = n2785 & n2804;
  assign n2806 = ~x591 & ~x592;
  assign n2807 = ~n2805 & n2806;
  assign n2808 = ~n2766 & ~n2807;
  assign n2809 = ~x591 & n2703;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = n2810 ^ x588;
  assign n2812 = n2811 ^ x588;
  assign n2818 = x421 ^ x420;
  assign n2819 = n2818 ^ x419;
  assign n2816 = x459 ^ x454;
  assign n2814 = x432 ^ x425;
  assign n2813 = x424 ^ x423;
  assign n2815 = n2814 ^ n2813;
  assign n2817 = n2816 ^ n2815;
  assign n2820 = n2819 ^ n2817;
  assign n2821 = x1198 & n2820;
  assign n2827 = x417 ^ x416;
  assign n2828 = n2827 ^ x415;
  assign n2825 = x464 ^ x453;
  assign n2823 = x431 ^ x418;
  assign n2822 = x438 ^ x437;
  assign n2824 = n2823 ^ n2822;
  assign n2826 = n2825 ^ n2824;
  assign n2829 = n2828 ^ n2826;
  assign n2830 = x1197 & n2829;
  assign n2831 = ~n2821 & ~n2830;
  assign n2837 = x428 ^ x427;
  assign n2838 = n2837 ^ x426;
  assign n2835 = x451 ^ x449;
  assign n2833 = x433 ^ x430;
  assign n2832 = x448 ^ x445;
  assign n2834 = n2833 ^ n2832;
  assign n2836 = n2835 ^ n2834;
  assign n2839 = n2838 ^ n2836;
  assign n2840 = x1199 & n2839;
  assign n2846 = x429 ^ x422;
  assign n2847 = n2846 ^ x414;
  assign n2844 = x443 ^ x436;
  assign n2842 = x446 ^ x444;
  assign n2841 = x435 ^ x434;
  assign n2843 = n2842 ^ n2841;
  assign n2845 = n2844 ^ n2843;
  assign n2848 = n2847 ^ n2845;
  assign n2849 = x1196 & n2848;
  assign n2850 = ~n2840 & ~n2849;
  assign n2851 = n2831 & n2850;
  assign n2852 = x588 & n2703;
  assign n2853 = ~n2851 & n2852;
  assign n2854 = n2853 ^ x588;
  assign n2855 = ~n2812 & ~n2854;
  assign n2856 = n2855 ^ x588;
  assign n2857 = ~x217 & ~n2856;
  assign n2858 = ~n2725 & n2857;
  assign n2859 = n1474 & n2858;
  assign n2860 = ~n2681 & ~n2859;
  assign n2861 = ~n2642 & n2860;
  assign n2862 = ~n2702 & n2857;
  assign n2863 = ~x286 & ~x289;
  assign n2864 = ~x285 & ~x288;
  assign n2865 = n2863 & n2864;
  assign n2866 = ~n2862 & ~n2865;
  assign n2867 = ~n2861 & ~n2866;
  assign n2868 = x1092 & x1093;
  assign n2869 = ~x98 & x567;
  assign n2870 = n2868 & ~n2869;
  assign n2871 = ~x1161 & ~x1162;
  assign n2872 = ~x1163 & n2871;
  assign n2873 = ~n2870 & n2872;
  assign n2874 = n1571 & n2873;
  assign n2875 = ~n2867 & n2874;
  assign n2876 = x567 & n2320;
  assign n2877 = ~x1199 & ~n2876;
  assign n2878 = ~x217 & ~x588;
  assign n2879 = x591 & ~x1091;
  assign n2880 = n2878 & n2879;
  assign n2881 = ~n2877 & n2880;
  assign n2882 = n2700 & n2881;
  assign n2883 = n2723 & n2882;
  assign n2884 = n1474 & n2317;
  assign n2885 = n2635 & n2884;
  assign n2886 = n2885 ^ n2639;
  assign n2887 = n2609 & n2886;
  assign n2888 = n2887 ^ n2639;
  assign n2889 = ~n2883 & n2888;
  assign n2890 = ~n2633 & ~n2889;
  assign n2891 = ~n2680 & ~n2890;
  assign n2892 = ~n1584 & ~n2390;
  assign n2893 = n2661 & n2892;
  assign n2894 = ~x122 & n2884;
  assign n2895 = ~x98 & n2894;
  assign n2896 = ~n2893 & ~n2895;
  assign n2897 = n2876 & n2883;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = ~n2891 & ~n2898;
  assign n2900 = n2875 & ~n2899;
  assign n2901 = ~n2865 & n2894;
  assign n2902 = n2869 & n2871;
  assign n2903 = n2901 & n2902;
  assign n2904 = ~n1571 & n2903;
  assign n2905 = ~n2858 & n2904;
  assign n2906 = ~x31 & n2868;
  assign n2907 = x1161 & x1162;
  assign n2908 = n2906 & n2907;
  assign n2909 = ~n2905 & ~n2908;
  assign n2910 = ~x1163 & ~n2909;
  assign n2911 = ~n2900 & ~n2910;
  assign n2912 = x76 & n1395;
  assign n2913 = ~n1478 & ~n2865;
  assign n2914 = ~x137 & ~n1259;
  assign n2915 = ~x50 & n2914;
  assign n2916 = ~n2913 & n2915;
  assign n2917 = n2912 & n2916;
  assign n2918 = ~x24 & n1233;
  assign n2919 = x50 & n2918;
  assign n2920 = ~x841 & n1259;
  assign n2921 = x32 & ~x841;
  assign n2922 = ~x24 & n2921;
  assign n2923 = n2922 ^ x32;
  assign n2924 = ~n2920 & n2923;
  assign n2925 = ~n2919 & ~n2924;
  assign n2926 = ~n2917 & n2925;
  assign n2927 = n1752 & ~n2926;
  assign n2928 = ~x252 & n1496;
  assign n2929 = n2320 ^ x129;
  assign n2930 = n2316 & n2929;
  assign n2931 = n2930 ^ x129;
  assign n2932 = n2473 & n2931;
  assign n2933 = ~n2928 & n2932;
  assign n2934 = x252 & ~n2650;
  assign n2935 = x75 & n2652;
  assign n2936 = ~n1478 & n2935;
  assign n2937 = ~n2934 & n2936;
  assign n2938 = ~n2933 & ~n2937;
  assign n2939 = n1496 & n2936;
  assign n2940 = n2650 & ~n2939;
  assign n2941 = ~x137 & ~n2940;
  assign n2942 = ~n2938 & n2941;
  assign n2943 = n2472 & n2942;
  assign n2944 = ~n2927 & ~n2943;
  assign n2945 = ~x70 & n1287;
  assign n2946 = ~n1455 & ~n2945;
  assign n2947 = n1326 & ~n2449;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = x73 & n2439;
  assign n2950 = n1253 & n1264;
  assign n2951 = n2949 & n2950;
  assign n2952 = n2948 & ~n2951;
  assign n2953 = ~x195 & ~x196;
  assign n2954 = ~x138 & ~x139;
  assign n2955 = n2953 & n2954;
  assign n2956 = ~x79 & ~x118;
  assign n2957 = ~x33 & ~x34;
  assign n2958 = n2956 & n2957;
  assign n2959 = n2955 & n2958;
  assign n2960 = x954 ^ x33;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = ~x63 & ~x107;
  assign n2963 = ~x40 & n2962;
  assign n2964 = ~n2961 & n2963;
  assign n2965 = x186 ^ x164;
  assign n2966 = ~x299 & n2965;
  assign n2967 = n2966 ^ x164;
  assign n2968 = n2643 & n2967;
  assign n2969 = ~n1563 & ~n2968;
  assign n2970 = n1593 & ~n2969;
  assign n2971 = n2964 & n2970;
  assign n2972 = n2952 & n2971;
  assign n2973 = n1264 & n2441;
  assign n2974 = ~n2385 & ~n2481;
  assign n2975 = ~n2379 & ~n2974;
  assign n2976 = n2973 & n2975;
  assign n2977 = n1565 & n2976;
  assign n2978 = x39 & n2643;
  assign n2979 = n2643 ^ n1574;
  assign n2980 = ~n2360 & n2364;
  assign n2981 = ~x174 & n2980;
  assign n2982 = n2367 & ~n2374;
  assign n2983 = ~x152 & n2982;
  assign n2984 = ~n2981 & ~n2983;
  assign n2985 = n2481 & ~n2984;
  assign n2986 = x176 & n2980;
  assign n2987 = x154 & n2982;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = n2385 & ~n2988;
  assign n2990 = ~n2985 & ~n2989;
  assign n2991 = n2990 ^ n2978;
  assign n2992 = n2979 & n2991;
  assign n2993 = n2992 ^ n2990;
  assign n2994 = n2978 & n2993;
  assign n2995 = n2994 ^ n2643;
  assign n2996 = n2977 & ~n2995;
  assign n2997 = n1589 & n2973;
  assign n2998 = ~n1566 & n2964;
  assign n2999 = n2998 ^ x92;
  assign n3000 = n2999 ^ n2998;
  assign n3001 = x176 ^ x154;
  assign n3002 = ~x299 & n3001;
  assign n3003 = n3002 ^ x154;
  assign n3004 = n2643 & n3003;
  assign n3005 = n2963 & n3004;
  assign n3006 = n3005 ^ n2998;
  assign n3007 = n3006 ^ n2998;
  assign n3008 = n3000 & n3007;
  assign n3009 = n3008 ^ n2998;
  assign n3010 = n2997 & n3009;
  assign n3011 = n3010 ^ n2998;
  assign n3012 = ~n2996 & n3011;
  assign n3013 = n1565 & n2635;
  assign n3014 = n2627 & n3013;
  assign n3015 = x38 & ~n3014;
  assign n3016 = ~x54 & ~n3015;
  assign n3017 = ~n3012 & n3016;
  assign n3018 = ~x74 & ~n2969;
  assign n3019 = ~n3017 & n3018;
  assign n3020 = x191 ^ x169;
  assign n3021 = ~x299 & n3020;
  assign n3022 = n3021 ^ x169;
  assign n3023 = n2643 & n3022;
  assign n3024 = x74 & n3023;
  assign n3025 = n1561 & ~n3024;
  assign n3026 = ~n3019 & n3025;
  assign n3027 = ~n1561 & n2643;
  assign n3029 = x183 ^ x178;
  assign n3028 = x157 ^ x149;
  assign n3030 = n3029 ^ n3028;
  assign n3031 = ~x299 & n3030;
  assign n3032 = n3031 ^ n3028;
  assign n3033 = n3027 & n3032;
  assign n3034 = ~n3026 & ~n3033;
  assign n3035 = n1571 & ~n3034;
  assign n3036 = ~n2972 & n3035;
  assign n3037 = n1326 & n2447;
  assign n3038 = x193 ^ x172;
  assign n3039 = ~x299 & n3038;
  assign n3040 = n3039 ^ x172;
  assign n3041 = n3037 & n3040;
  assign n3042 = x180 ^ x158;
  assign n3043 = ~x299 & n3042;
  assign n3044 = n3043 ^ x158;
  assign n3045 = n1284 & n3044;
  assign n3046 = n1254 & n3045;
  assign n3047 = ~x198 & ~x299;
  assign n3048 = ~x841 & n1205;
  assign n3049 = n3047 & n3048;
  assign n3050 = n2441 & n3049;
  assign n3051 = ~x299 & ~n2945;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = x183 & ~n3052;
  assign n3057 = x299 ^ x152;
  assign n3058 = n3057 ^ x152;
  assign n3059 = x174 ^ x152;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = n3060 ^ x152;
  assign n3062 = n3061 ^ x299;
  assign n3054 = ~x210 & n2921;
  assign n3055 = n2945 & ~n3054;
  assign n3056 = x149 & ~n3055;
  assign n3063 = n3062 ^ n3056;
  assign n3064 = n3063 ^ n3062;
  assign n3065 = n3062 ^ n3061;
  assign n3066 = n3064 & n3065;
  assign n3067 = n3066 ^ n3062;
  assign n3068 = ~x73 & n3067;
  assign n3069 = n3068 ^ n3062;
  assign n3070 = ~n3053 & ~n3069;
  assign n3071 = ~n3046 & n3070;
  assign n3072 = ~n3041 & n3071;
  assign n3073 = ~n1463 & ~n3072;
  assign n3074 = ~x39 & ~n3073;
  assign n3075 = n1658 & n2995;
  assign n3076 = ~n3074 & n3075;
  assign n3077 = n3036 & ~n3076;
  assign n3078 = n1563 & n1570;
  assign n3079 = n1562 & n3078;
  assign n3080 = n2963 & n3079;
  assign n3081 = n1568 & n1575;
  assign n3082 = x149 & n2643;
  assign n3083 = n3082 ^ n2961;
  assign n3084 = n3081 & ~n3083;
  assign n3085 = n3084 ^ n2961;
  assign n3086 = n3080 & ~n3085;
  assign n3087 = n3028 ^ n1561;
  assign n3088 = n3087 ^ n3028;
  assign n3089 = n3078 ^ x169;
  assign n3090 = n3089 ^ x169;
  assign n3091 = x169 ^ x164;
  assign n3092 = n3091 ^ x169;
  assign n3093 = ~n3090 & n3092;
  assign n3094 = n3093 ^ x169;
  assign n3095 = ~x74 & n3094;
  assign n3096 = n3095 ^ x169;
  assign n3097 = n3096 ^ n3028;
  assign n3098 = n3088 & n3097;
  assign n3099 = n3098 ^ n3028;
  assign n3100 = n2643 & n3099;
  assign n3101 = n3100 ^ n1561;
  assign n3102 = ~n1571 & n3101;
  assign n3103 = ~n3086 & n3102;
  assign n3104 = ~n3077 & ~n3103;
  assign n3105 = n1572 & n2952;
  assign n3106 = n1566 & n1568;
  assign n3107 = n2973 & n3106;
  assign n3108 = ~n1569 & ~n3107;
  assign n3109 = ~n3105 & ~n3108;
  assign n3110 = ~x33 & ~x954;
  assign n3111 = n3110 ^ x34;
  assign n3112 = n2959 & n3110;
  assign n3113 = n3111 & n3112;
  assign n3114 = n3113 ^ n3111;
  assign n3115 = ~n3109 & ~n3114;
  assign n3116 = ~x144 & n2980;
  assign n3117 = ~x161 & n2982;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = n2480 & ~n3118;
  assign n3120 = x177 & n2980;
  assign n3121 = x155 & n2982;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = n1481 & ~n3122;
  assign n3124 = ~n3119 & ~n3123;
  assign n3125 = n2643 & ~n3124;
  assign n3126 = n2977 & ~n3125;
  assign n3127 = ~n1567 & n1569;
  assign n3128 = ~n3126 & n3127;
  assign n3129 = x39 & n2977;
  assign n3130 = x92 & n2997;
  assign n3131 = n3130 ^ n3114;
  assign n3132 = n3131 ^ n3114;
  assign n3133 = x177 ^ x155;
  assign n3134 = ~x299 & n3133;
  assign n3135 = n3134 ^ x155;
  assign n3136 = n2643 & n3135;
  assign n3137 = n3136 ^ n3114;
  assign n3138 = n3132 & ~n3137;
  assign n3139 = n3138 ^ n3114;
  assign n3140 = ~n3129 & n3139;
  assign n3141 = n3128 & ~n3140;
  assign n3142 = ~n3115 & ~n3141;
  assign n3143 = n3080 & ~n3142;
  assign n3144 = ~n1490 & ~n1494;
  assign n3145 = n3037 & ~n3144;
  assign n3146 = x140 & ~n3052;
  assign n3147 = x162 & x299;
  assign n3148 = ~n3055 & n3147;
  assign n3149 = x181 ^ x159;
  assign n3150 = ~x299 & n3149;
  assign n3151 = n3150 ^ x159;
  assign n3152 = n2442 & n3151;
  assign n3153 = x299 ^ x144;
  assign n3154 = n3153 ^ x144;
  assign n3155 = x161 ^ x144;
  assign n3156 = n3154 & n3155;
  assign n3157 = n3156 ^ x144;
  assign n3158 = x73 & ~n3157;
  assign n3159 = ~n3152 & ~n3158;
  assign n3160 = ~n3148 & n3159;
  assign n3161 = ~n3146 & n3160;
  assign n3162 = ~n3145 & n3161;
  assign n3163 = n1752 & ~n3162;
  assign n3176 = x197 ^ x162;
  assign n3175 = ~x149 & ~x157;
  assign n3177 = n3176 ^ n3175;
  assign n3178 = n3177 ^ n1729;
  assign n3179 = n3178 ^ n3177;
  assign n3181 = x145 ^ x140;
  assign n3180 = ~x178 & ~x183;
  assign n3182 = n3181 ^ n3180;
  assign n3183 = n3182 ^ n3177;
  assign n3184 = n3179 & n3183;
  assign n3185 = n3184 ^ n3177;
  assign n3164 = x188 ^ x167;
  assign n3165 = ~x299 & n3164;
  assign n3166 = n3165 ^ x167;
  assign n3167 = ~x74 & n3166;
  assign n3168 = ~n3016 & n3167;
  assign n3169 = x148 ^ x141;
  assign n3170 = x299 & n3169;
  assign n3171 = n3170 ^ x141;
  assign n3172 = x74 & n3171;
  assign n3173 = n1571 & ~n3172;
  assign n3174 = ~n3168 & n3173;
  assign n3186 = n3185 ^ n3174;
  assign n3187 = n3186 ^ n3185;
  assign n3188 = ~x74 & ~n3078;
  assign n3189 = x167 & n3188;
  assign n3190 = x74 & x148;
  assign n3191 = ~n1571 & ~n3190;
  assign n3192 = ~n3189 & n3191;
  assign n3193 = n3192 ^ n3185;
  assign n3194 = n3193 ^ n3185;
  assign n3195 = ~n3187 & ~n3194;
  assign n3196 = n3195 ^ n3185;
  assign n3197 = n1561 & ~n3196;
  assign n3198 = n3197 ^ n3185;
  assign n3199 = ~n3163 & n3198;
  assign n3200 = n1633 & n3107;
  assign n3201 = x162 & n3200;
  assign n3202 = n3199 & ~n3201;
  assign n3203 = n2643 & ~n3202;
  assign n3204 = ~n3143 & ~n3203;
  assign n3205 = x24 & x59;
  assign n3206 = ~x55 & ~x74;
  assign n3207 = ~n3205 & n3206;
  assign n3208 = n1596 & n3207;
  assign n3209 = x841 ^ x93;
  assign n3210 = n1451 & n3209;
  assign n3211 = n2428 & ~n3210;
  assign n3212 = ~x122 & n2320;
  assign n3213 = ~n2913 & n3212;
  assign n3214 = x76 & ~n2914;
  assign n3215 = n3213 & n3214;
  assign n3216 = ~n1503 & ~n3215;
  assign n3217 = ~n3211 & ~n3216;
  assign n3218 = x40 & x1082;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = ~n1463 & ~n3219;
  assign n3221 = n1597 & ~n2436;
  assign n3222 = x24 & ~x59;
  assign n3223 = ~n3221 & ~n3222;
  assign n3224 = ~n3220 & ~n3223;
  assign n3229 = ~n1496 & ~n2331;
  assign n3227 = x137 & ~n1478;
  assign n3228 = ~n2934 & ~n3227;
  assign n3230 = n3229 ^ n3228;
  assign n3231 = x75 ^ x38;
  assign n3232 = n3231 ^ n3229;
  assign n3233 = ~n3229 & ~n3232;
  assign n3234 = n3233 ^ n3229;
  assign n3235 = n3230 & ~n3234;
  assign n3236 = n3235 ^ n3233;
  assign n3237 = n3236 ^ n3229;
  assign n3238 = n3237 ^ n3231;
  assign n3239 = x75 & ~n3238;
  assign n3240 = n3239 ^ n3231;
  assign n3241 = n2652 & n3240;
  assign n3242 = n2389 & n2650;
  assign n3243 = x683 & n3242;
  assign n3244 = x137 & n2934;
  assign n3245 = n3244 ^ x252;
  assign n3246 = ~n3243 & n3245;
  assign n3247 = ~x137 & ~n1496;
  assign n3248 = n1563 & ~n3247;
  assign n3249 = ~n3229 & n3248;
  assign n3250 = n2932 & n3249;
  assign n3251 = ~n3246 & n3250;
  assign n3252 = ~n3241 & ~n3251;
  assign n3253 = n3014 & ~n3252;
  assign n3225 = ~n3014 & n3188;
  assign n3226 = n1592 & ~n3225;
  assign n3254 = n3253 ^ n3226;
  assign n3255 = n3224 & n3254;
  assign n3256 = n3255 ^ n3226;
  assign n3257 = n3208 & n3256;
  assign n3258 = x36 & n1246;
  assign n3259 = n1395 & n3258;
  assign n3260 = ~n2619 & ~n3259;
  assign n3261 = n1252 & n2412;
  assign n3262 = ~n3260 & n3261;
  assign n3263 = ~n2320 & n3262;
  assign n3264 = n1246 & n3261;
  assign n3265 = n1395 & n3264;
  assign n3266 = ~x841 & n3265;
  assign n3267 = ~x70 & ~x89;
  assign n3268 = x332 & ~n3267;
  assign n3269 = n3266 & n3268;
  assign n3270 = n1431 & n3264;
  assign n3271 = x64 & n3270;
  assign n3272 = ~x841 & n3271;
  assign n3273 = ~n3269 & ~n3272;
  assign n3274 = x24 & n1588;
  assign n3275 = n3273 & ~n3274;
  assign n3276 = ~x35 & ~x48;
  assign n3277 = x841 ^ x47;
  assign n3278 = n3277 ^ x841;
  assign n3279 = ~x986 & n2320;
  assign n3280 = x252 & ~n3279;
  assign n3281 = x108 & x314;
  assign n3282 = ~n3280 & n3281;
  assign n3283 = n3282 ^ x841;
  assign n3284 = n3283 ^ x841;
  assign n3285 = ~n3278 & ~n3284;
  assign n3286 = n3285 ^ x841;
  assign n3287 = n3276 & n3286;
  assign n3288 = n3287 ^ x841;
  assign n3289 = n2435 & ~n3288;
  assign n3290 = n1256 & n2920;
  assign n3291 = n1572 & n3290;
  assign n3292 = ~x287 & n2567;
  assign n3293 = x835 & x984;
  assign n3294 = ~x979 & ~n3293;
  assign n3295 = ~n2382 & n3294;
  assign n3297 = x835 & ~n2396;
  assign n3298 = n2391 & n3297;
  assign n3296 = ~x1093 & ~n2394;
  assign n3299 = n3298 ^ n3296;
  assign n3300 = n3299 ^ n3296;
  assign n3301 = x786 & ~x1082;
  assign n3302 = n3295 & n3301;
  assign n3303 = n3302 ^ n3296;
  assign n3304 = ~n3300 & ~n3303;
  assign n3305 = n3304 ^ n3296;
  assign n3306 = n3295 & n3305;
  assign n3307 = n3292 & n3306;
  assign n3308 = ~n3291 & ~n3307;
  assign n3309 = ~n3289 & n3308;
  assign n3310 = x102 ^ x40;
  assign n3311 = ~x102 & x1082;
  assign n3312 = n3310 & n3311;
  assign n3313 = n3312 ^ n3310;
  assign n3314 = n1752 & n3313;
  assign n3315 = ~n1248 & ~n1478;
  assign n3316 = ~n2611 & ~n3315;
  assign n3317 = n2473 & ~n2673;
  assign n3318 = ~n1584 & ~n3317;
  assign n3319 = x228 & ~n3318;
  assign n3320 = ~n2625 & n3319;
  assign n3321 = ~n3316 & n3320;
  assign n3322 = x110 ^ x94;
  assign n3323 = ~x250 & x252;
  assign n3324 = x901 & ~x959;
  assign n3325 = n3323 & n3324;
  assign n3326 = n3325 ^ x110;
  assign n3327 = n3326 ^ n3325;
  assign n3328 = ~x480 & x949;
  assign n3329 = n3328 ^ n3325;
  assign n3330 = n3327 & n3329;
  assign n3331 = n3330 ^ n3325;
  assign n3332 = n3322 & n3331;
  assign n3333 = ~n2599 & n3332;
  assign n3334 = ~x87 & ~x100;
  assign n3335 = ~n1574 & ~n3334;
  assign n3336 = ~x228 & ~n3332;
  assign n3337 = x87 & x100;
  assign n3338 = n1657 & ~n3337;
  assign n3339 = n1571 & n3338;
  assign n3340 = ~n3336 & n3339;
  assign n3341 = ~n3335 & n3340;
  assign n3342 = ~n2657 & n3341;
  assign n3343 = ~n2632 & n3342;
  assign n3344 = ~n3333 & n3343;
  assign n3345 = ~n3321 & n3344;
  assign n3346 = ~x44 & n3345;
  assign n3347 = ~x101 & n3346;
  assign n3348 = n3347 ^ x41;
  assign n3349 = n2634 & ~n3348;
  assign n3350 = x287 & n2566;
  assign n3351 = n2562 & n3350;
  assign n3352 = n2643 & ~n3351;
  assign n3353 = n2563 & n3352;
  assign n3354 = x161 & ~n1729;
  assign n3355 = n1492 & n3354;
  assign n3356 = n3355 ^ n3352;
  assign n3357 = x144 & n1729;
  assign n3358 = n1488 & n3357;
  assign n3359 = n3358 ^ n3353;
  assign n3360 = ~n3356 & n3359;
  assign n3361 = n3360 ^ n3358;
  assign n3362 = n3353 & n3361;
  assign n3363 = n3362 ^ n2563;
  assign n3364 = ~n3349 & ~n3363;
  assign n3365 = n2324 & n3346;
  assign n3366 = n2328 & n3365;
  assign n3367 = ~x114 & n3366;
  assign n3368 = n3367 ^ x42;
  assign n3369 = n2634 & n3368;
  assign n3370 = ~x189 & n1729;
  assign n3371 = n3370 ^ n3352;
  assign n3372 = ~x166 & ~n1729;
  assign n3373 = n3372 ^ n3353;
  assign n3374 = ~n3371 & n3373;
  assign n3375 = n3374 ^ n3372;
  assign n3376 = n3353 & n3375;
  assign n3377 = n3376 ^ n2563;
  assign n3378 = ~x199 & ~x200;
  assign n3379 = ~x299 & ~n3378;
  assign n3380 = n1571 & n3379;
  assign n3381 = x207 & x208;
  assign n3382 = ~x199 & ~n3381;
  assign n3383 = n3380 & ~n3382;
  assign n3384 = x212 & x214;
  assign n3385 = x211 & n3384;
  assign n3386 = n3385 ^ x219;
  assign n3387 = n3385 ^ n1729;
  assign n3388 = ~n3385 & n3387;
  assign n3389 = n3388 ^ n3385;
  assign n3390 = n3386 & ~n3389;
  assign n3391 = n3390 ^ n3388;
  assign n3392 = n3391 ^ n3385;
  assign n3393 = n3392 ^ n1729;
  assign n3394 = ~n3383 & n3393;
  assign n3395 = n3394 ^ n3383;
  assign n3396 = n3377 & n3395;
  assign n3397 = ~n3369 & ~n3396;
  assign n3398 = ~x42 & n3367;
  assign n3399 = n3398 ^ x43;
  assign n3400 = n2634 & n3399;
  assign n3404 = ~x211 & ~x219;
  assign n3405 = n3404 ^ x211;
  assign n3406 = n3384 & n3405;
  assign n3407 = n3406 ^ x211;
  assign n3401 = n3378 ^ x200;
  assign n3402 = n3381 & n3401;
  assign n3403 = n3402 ^ x200;
  assign n3408 = n3407 ^ n3403;
  assign n3409 = ~n1729 & n3408;
  assign n3410 = n3409 ^ n3403;
  assign n3411 = n3377 & n3410;
  assign n3412 = ~n3400 & ~n3411;
  assign n3413 = n3345 ^ x44;
  assign n3414 = n2634 & n3413;
  assign n3415 = n1489 & n1729;
  assign n3416 = n1493 & ~n1729;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = n3353 & ~n3417;
  assign n3419 = ~n3414 & ~n3418;
  assign n3420 = x979 & n3292;
  assign n3421 = x46 & ~x109;
  assign n3422 = n2412 & n3421;
  assign n3423 = n1292 & n3422;
  assign n3424 = n1326 & n3423;
  assign n3425 = x24 & n3424;
  assign n3426 = x61 & n3266;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = ~n3265 & ~n3270;
  assign n3429 = ~x36 & ~x88;
  assign n3430 = ~x104 & n3429;
  assign n3431 = ~n2389 & ~n3430;
  assign n3432 = ~n3428 & n3431;
  assign n3433 = n3432 ^ n3261;
  assign n3434 = n3433 ^ n3432;
  assign n3435 = ~n1478 & ~n2318;
  assign n3436 = n3435 ^ n3432;
  assign n3437 = n3436 ^ n3432;
  assign n3438 = n3434 & n3437;
  assign n3439 = n3438 ^ n3432;
  assign n3440 = ~n3260 & n3439;
  assign n3441 = n3440 ^ n3432;
  assign n3442 = x841 & n3265;
  assign n3443 = x48 & n3442;
  assign n3444 = x74 & n2652;
  assign n3445 = n1613 & n3444;
  assign n3446 = x49 & n3442;
  assign n3447 = ~n3445 & ~n3446;
  assign n3448 = n1449 & n3261;
  assign n3449 = x24 & x50;
  assign n3450 = n3448 & n3449;
  assign n3451 = ~n2474 & ~n2936;
  assign n3452 = n3229 & ~n3451;
  assign n3453 = n2472 & n3452;
  assign n3454 = x94 & ~x110;
  assign n3455 = ~x58 & n3261;
  assign n3456 = ~x86 & n1236;
  assign n3457 = n1289 & n3456;
  assign n3458 = n3455 & n3457;
  assign n3459 = n1233 & n3458;
  assign n3460 = n3454 & n3459;
  assign n3461 = n2650 ^ n1478;
  assign n3462 = ~x252 & n3461;
  assign n3463 = n3462 ^ n1478;
  assign n3464 = n3460 & n3463;
  assign n3465 = ~n3453 & ~n3464;
  assign n3466 = ~n3450 & n3465;
  assign n3467 = n1334 & n1351;
  assign n3468 = n1393 & n3264;
  assign n3469 = n3467 & n3468;
  assign n3470 = x82 & ~x111;
  assign n3471 = n3469 & n3470;
  assign n3472 = n2330 & n3345;
  assign n3473 = n3472 ^ x52;
  assign n3474 = n2634 & n3473;
  assign n3475 = ~x211 & x219;
  assign n3476 = ~n1729 & ~n3475;
  assign n3477 = ~x219 & n3407;
  assign n3478 = x211 & ~x219;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = n3476 & n3479;
  assign n3481 = ~x199 & x200;
  assign n3482 = ~x299 & ~n3481;
  assign n3483 = n1571 & n3482;
  assign n3484 = ~x200 & ~n3382;
  assign n3485 = n3483 & ~n3484;
  assign n3486 = ~n3480 & ~n3485;
  assign n3487 = ~n3395 & ~n3486;
  assign n3488 = n3377 & n3487;
  assign n3489 = ~n3474 & ~n3488;
  assign n3490 = ~x979 & n3293;
  assign n3491 = n3292 & n3490;
  assign n3492 = n1240 & n3455;
  assign n3493 = n2297 & n3492;
  assign n3494 = x53 & ~x60;
  assign n3495 = n3493 & n3494;
  assign n3496 = x24 & n3495;
  assign n3497 = ~n3491 & ~n3496;
  assign n3498 = x24 & n1614;
  assign n3499 = n1593 & n3498;
  assign n3500 = x106 & n3266;
  assign n3501 = ~n3499 & ~n3500;
  assign n3502 = x24 & n3200;
  assign n3503 = x45 & n3265;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = ~x62 & x841;
  assign n3506 = n1617 & n3505;
  assign n3507 = x55 & ~x56;
  assign n3508 = ~x24 & ~x62;
  assign n3509 = n3507 & n3508;
  assign n3510 = ~n3506 & ~n3509;
  assign n3511 = n1576 & ~n3510;
  assign n3512 = ~x841 & n1618;
  assign n3513 = x62 & x924;
  assign n3514 = n3512 & ~n3513;
  assign n3515 = x24 & n1580;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = n1247 & n2413;
  assign n3518 = ~x841 & n3517;
  assign n3519 = n3512 & n3513;
  assign n3520 = ~x57 & n1569;
  assign n3521 = n3205 & n3520;
  assign n3522 = n1575 & n3521;
  assign n3523 = ~n3519 & ~n3522;
  assign n3524 = n2382 & n3294;
  assign n3525 = n3292 & n3524;
  assign n3526 = ~x53 & x60;
  assign n3527 = n3493 & n3526;
  assign n3528 = x24 & n3527;
  assign n3529 = ~n3525 & ~n3528;
  assign n3530 = x61 & n3442;
  assign n3531 = ~x24 & n3527;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = x62 & x841;
  assign n3534 = n3533 ^ n3508;
  assign n3535 = ~x57 & n3534;
  assign n3536 = n3535 ^ n3508;
  assign n3537 = ~n1632 & n3536;
  assign n3538 = ~x24 & n3424;
  assign n3539 = x63 & n3270;
  assign n3540 = x999 & n3539;
  assign n3541 = ~n3538 & ~n3540;
  assign n3542 = x841 & n3271;
  assign n3543 = x107 & n3270;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = ~n3298 & n3302;
  assign n3546 = n3292 & n3545;
  assign n3547 = n1396 & n3264;
  assign n3548 = x81 & n1224;
  assign n3549 = x314 & n1226;
  assign n3550 = n3548 & n3549;
  assign n3551 = n3547 & n3550;
  assign n3552 = x219 ^ x199;
  assign n3553 = x299 & n3552;
  assign n3554 = n3553 ^ x199;
  assign n3555 = n3551 & n3554;
  assign n3556 = ~x69 & n1384;
  assign n3557 = n3468 & n3556;
  assign n3558 = x314 & n3557;
  assign n3559 = x83 & ~x103;
  assign n3560 = n3558 & n3559;
  assign n3561 = n2481 & n2567;
  assign n3562 = n1779 & ~n2363;
  assign n3563 = x299 & n1741;
  assign n3564 = ~n2377 & n3563;
  assign n3565 = ~n3562 & ~n3564;
  assign n3566 = n3561 & ~n3565;
  assign n3567 = x69 & ~x314;
  assign n3568 = ~x71 & ~n3567;
  assign n3569 = n3265 & ~n3568;
  assign n3570 = x24 & x70;
  assign n3571 = n2435 & n3570;
  assign n3572 = n2385 & n2567;
  assign n3573 = ~n3561 & ~n3572;
  assign n3574 = n1534 & ~n2377;
  assign n3575 = x210 & n3574;
  assign n3576 = n1538 & ~n2363;
  assign n3577 = x198 & n3576;
  assign n3578 = ~n3575 & ~n3577;
  assign n3579 = x589 & ~n3578;
  assign n3580 = ~n3573 & n3579;
  assign n3581 = ~x593 & n3580;
  assign n3582 = n2564 & n3350;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = ~n3571 & n3583;
  assign n3585 = n3481 ^ n3478;
  assign n3586 = ~x299 & n3585;
  assign n3587 = n3586 ^ n3478;
  assign n3588 = n3551 & n3587;
  assign n3589 = ~n1354 & n3468;
  assign n3590 = x85 & n1332;
  assign n3591 = n1369 & n3590;
  assign n3592 = ~n1362 & n3591;
  assign n3593 = x314 & n3592;
  assign n3594 = n3589 & n3593;
  assign n3595 = ~n3588 & ~n3594;
  assign n3596 = x88 & n2477;
  assign n3597 = ~n1455 & n3596;
  assign n3598 = ~x38 & ~n3597;
  assign n3599 = x72 & n1282;
  assign n3600 = x24 & n3599;
  assign n3601 = n3598 & ~n3600;
  assign n3602 = n1572 & ~n3601;
  assign n3603 = n2670 & n3561;
  assign n3604 = ~n3602 & ~n3603;
  assign n3605 = x73 & n1752;
  assign n3606 = ~n2379 & n3561;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~x314 & x1050;
  assign n3609 = ~x39 & ~n3608;
  assign n3610 = ~n3607 & ~n3609;
  assign n3611 = x479 & n1259;
  assign n3612 = n2320 & ~n3611;
  assign n3613 = ~x96 & ~n3612;
  assign n3614 = ~x479 & ~x841;
  assign n3615 = x96 & ~n3614;
  assign n3616 = ~n1478 & ~n3615;
  assign n3617 = n1572 & n3616;
  assign n3618 = ~n3613 & n3617;
  assign n3619 = ~n1470 & n3618;
  assign n3620 = x74 & n3498;
  assign n3621 = ~n3619 & ~n3620;
  assign n3622 = n1487 & n1572;
  assign n3623 = x75 & n3498;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = n2865 & n2914;
  assign n3626 = ~n3213 & ~n3625;
  assign n3627 = n2912 & n3626;
  assign n3628 = x94 & ~n2650;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = x252 ^ x94;
  assign n3631 = n3630 ^ x252;
  assign n3632 = n2914 ^ x252;
  assign n3633 = ~n3631 & n3632;
  assign n3634 = n3633 ^ x252;
  assign n3635 = n1478 & n3634;
  assign n3636 = ~n3629 & ~n3635;
  assign n3637 = n1752 & n3636;
  assign n3638 = x77 & x314;
  assign n3639 = ~n1237 & ~n3638;
  assign n3640 = n2435 & n3639;
  assign n3641 = x232 & n2590;
  assign n3645 = ~x166 & n2962;
  assign n3646 = n2949 & n3645;
  assign n3647 = ~x163 & x299;
  assign n3648 = ~n3646 & n3647;
  assign n3649 = ~n3037 & ~n3648;
  assign n3650 = x153 & n1305;
  assign n3651 = n2446 & n3650;
  assign n3652 = ~x40 & x95;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = n3653 ^ x175;
  assign n3655 = n3654 ^ x175;
  assign n3656 = n1503 ^ x175;
  assign n3657 = n3656 ^ x175;
  assign n3658 = ~n3655 & n3657;
  assign n3659 = n3658 ^ x175;
  assign n3660 = x299 & n3659;
  assign n3661 = n3660 ^ x175;
  assign n3662 = ~n3649 & ~n3661;
  assign n3663 = x189 ^ x166;
  assign n3664 = ~x299 & n3663;
  assign n3665 = n3664 ^ x166;
  assign n3666 = n2951 & n3665;
  assign n3667 = n2643 & ~n3666;
  assign n3668 = x182 ^ x160;
  assign n3669 = ~x299 & n3668;
  assign n3670 = n3669 ^ x160;
  assign n3671 = n2443 & ~n3670;
  assign n3672 = n3667 & ~n3671;
  assign n3673 = ~x184 & ~n3052;
  assign n3674 = n3672 & ~n3673;
  assign n3675 = ~n3662 & n3674;
  assign n3642 = ~x34 & n3110;
  assign n3643 = n3642 ^ x79;
  assign n3644 = ~n2959 & n3643;
  assign n3676 = n3675 ^ n3644;
  assign n3677 = ~n2952 & ~n3676;
  assign n3678 = n3677 ^ n3644;
  assign n3679 = ~x39 & n3678;
  assign n3680 = ~n2976 & ~n3644;
  assign n3681 = ~x189 & n2980;
  assign n3682 = ~x166 & n2982;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n2481 & ~n3683;
  assign n3685 = x179 & n2980;
  assign n3686 = x156 & n2982;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = n2385 & ~n3687;
  assign n3689 = ~n3684 & ~n3688;
  assign n3690 = n2643 & ~n3689;
  assign n3691 = n2973 & n3690;
  assign n3692 = x39 & ~n3691;
  assign n3693 = ~n3680 & n3692;
  assign n3694 = n1565 & n2962;
  assign n3695 = ~x38 & n3694;
  assign n3696 = ~n3693 & n3695;
  assign n3697 = ~n3679 & n3696;
  assign n3698 = n3644 ^ n3130;
  assign n3699 = n3698 ^ n3644;
  assign n3700 = x179 ^ x156;
  assign n3701 = ~x299 & n3700;
  assign n3702 = n3701 ^ x156;
  assign n3703 = n2643 & n3702;
  assign n3704 = n3703 ^ n3644;
  assign n3705 = n3699 & ~n3704;
  assign n3706 = n3705 ^ n3644;
  assign n3707 = n2962 & ~n3706;
  assign n3708 = n1564 & ~n3707;
  assign n3709 = ~n1585 & ~n3708;
  assign n3710 = ~x40 & ~n3015;
  assign n3711 = ~n3709 & n3710;
  assign n3712 = ~n3697 & n3711;
  assign n3717 = n3180 ^ x145;
  assign n3718 = n3181 & n3717;
  assign n3719 = n3718 ^ x140;
  assign n3720 = n3719 ^ x184;
  assign n3713 = n3175 ^ x197;
  assign n3714 = n3176 & n3713;
  assign n3715 = n3714 ^ x162;
  assign n3716 = n3715 ^ x163;
  assign n3721 = n3720 ^ n3716;
  assign n3722 = ~x299 & n3721;
  assign n3723 = n3722 ^ n3716;
  assign n3724 = n3027 & n3723;
  assign n3725 = n1562 & ~n1563;
  assign n3726 = x187 ^ x147;
  assign n3727 = ~x299 & n3726;
  assign n3728 = n3727 ^ x147;
  assign n3729 = n2643 & n3728;
  assign n3730 = n3725 & ~n3729;
  assign n3731 = ~n3724 & ~n3730;
  assign n3732 = ~n3712 & n3731;
  assign n3733 = n1571 & ~n3732;
  assign n3734 = x163 & n2643;
  assign n3735 = n3734 ^ n3644;
  assign n3736 = n3107 & ~n3735;
  assign n3737 = n3736 ^ n3644;
  assign n3738 = n2962 & ~n3737;
  assign n3739 = ~x40 & ~n1569;
  assign n3740 = n3079 & n3739;
  assign n3741 = ~n3738 & n3740;
  assign n3742 = n3027 & n3716;
  assign n3743 = x147 & n2643;
  assign n3744 = n1562 & ~n3743;
  assign n3745 = ~n3742 & ~n3744;
  assign n3746 = ~n1571 & ~n3079;
  assign n3747 = ~n3745 & n3746;
  assign n3748 = ~n3741 & ~n3747;
  assign n3749 = ~n3733 & n3748;
  assign n3750 = ~x63 & ~n2414;
  assign n3751 = n1632 & ~n3750;
  assign n3752 = ~x592 & ~n2722;
  assign n3753 = n2702 & ~n3752;
  assign n3754 = ~x588 & ~x590;
  assign n3755 = n2700 & ~n3754;
  assign n3756 = x98 & ~x592;
  assign n3757 = x1199 & n3756;
  assign n3758 = n3757 ^ n2865;
  assign n3759 = n3757 ^ x590;
  assign n3760 = n3759 ^ x590;
  assign n3761 = n2894 ^ x590;
  assign n3762 = n3760 & ~n3761;
  assign n3763 = n3762 ^ x590;
  assign n3764 = n3758 & ~n3763;
  assign n3765 = n3764 ^ n2865;
  assign n3766 = ~n3755 & ~n3765;
  assign n3767 = n3753 & n3766;
  assign n3768 = n2561 & n2885;
  assign n3769 = ~n3767 & n3768;
  assign n3770 = ~n2637 & n3769;
  assign n3771 = ~n3751 & n3770;
  assign n3772 = n3753 & ~n3757;
  assign n3773 = n2901 & ~n3772;
  assign n3774 = ~n3771 & ~n3773;
  assign n3775 = n2857 & ~n3774;
  assign n3776 = ~n2870 & ~n3775;
  assign n3777 = ~x80 & n2872;
  assign n3778 = ~n3776 & n3777;
  assign n3779 = x81 & ~x314;
  assign n3780 = ~x68 & ~n3779;
  assign n3781 = ~n3428 & ~n3780;
  assign n3782 = x314 ^ x66;
  assign n3783 = x69 & n3782;
  assign n3784 = n3783 ^ x66;
  assign n3785 = n3265 & n3784;
  assign n3786 = ~x68 & x84;
  assign n3787 = n1229 & n3786;
  assign n3788 = n3589 & n3787;
  assign n3789 = ~x314 & n3559;
  assign n3790 = n3557 & n3789;
  assign n3791 = ~n3788 & ~n3790;
  assign n3792 = n3404 ^ n3378;
  assign n3793 = x299 & n3792;
  assign n3794 = n3793 ^ n3378;
  assign n3795 = n3551 & n3794;
  assign n3796 = ~x314 & n3592;
  assign n3797 = ~x67 & ~n3796;
  assign n3798 = n3589 & ~n3797;
  assign n3799 = ~n3565 & n3572;
  assign n3800 = n2426 & n3558;
  assign n3801 = x104 & n2389;
  assign n3802 = n3265 & n3801;
  assign n3803 = n2865 & n3802;
  assign n3804 = x88 & n2318;
  assign n3805 = n3270 & n3804;
  assign n3806 = ~n3803 & ~n3805;
  assign n3807 = x89 & x841;
  assign n3808 = ~x24 & x70;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = n2435 & ~n3809;
  assign n3811 = ~x1050 & n3605;
  assign n3812 = x841 & n3517;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = n2617 ^ n1481;
  assign n3815 = n2617 ^ x24;
  assign n3816 = n3815 ^ x24;
  assign n3817 = n3259 ^ x24;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = n3818 ^ x24;
  assign n3820 = n3814 & n3819;
  assign n3821 = n3820 ^ n1481;
  assign n3822 = n3455 & n3821;
  assign n3823 = n2567 & n2671;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = n3608 ^ n2386;
  assign n3826 = n3825 ^ n2386;
  assign n3827 = n2386 ^ x92;
  assign n3828 = n3827 ^ n2386;
  assign n3829 = n3826 & n3828;
  assign n3830 = n3829 ^ n2386;
  assign n3831 = ~x39 & n3830;
  assign n3832 = n3831 ^ n2386;
  assign n3833 = n1630 & n3832;
  assign n3834 = n2300 & n2435;
  assign n3835 = n1604 & n1653;
  assign n3836 = ~x1050 & n3835;
  assign n3837 = ~n3834 & ~n3836;
  assign n3838 = x49 & n3266;
  assign n3839 = ~n1478 & n2651;
  assign n3840 = n3460 & n3839;
  assign n3841 = ~n3838 & ~n3840;
  assign n3842 = ~n3574 & ~n3576;
  assign n3843 = ~n3573 & ~n3842;
  assign n3844 = ~n3579 & n3843;
  assign n3845 = x89 & ~x332;
  assign n3846 = n3266 & n3845;
  assign n3847 = ~n3844 & ~n3846;
  assign n3848 = ~x32 & ~x40;
  assign n3849 = n1572 & n3848;
  assign n3850 = x95 & n3849;
  assign n3851 = n1254 & n3850;
  assign n3852 = x24 & n3851;
  assign n3853 = n3847 & ~n3852;
  assign n3854 = ~n1254 & n1455;
  assign n3855 = x96 ^ x95;
  assign n3856 = x96 ^ x24;
  assign n3857 = n3856 ^ x24;
  assign n3858 = n3857 ^ n3855;
  assign n3859 = n3614 ^ n1479;
  assign n3860 = ~n1479 & n3859;
  assign n3861 = n3860 ^ x24;
  assign n3862 = n3861 ^ n1479;
  assign n3863 = n3858 & n3862;
  assign n3864 = n3863 ^ n3860;
  assign n3865 = n3864 ^ n1479;
  assign n3866 = n3855 & ~n3865;
  assign n3867 = n3849 & n3866;
  assign n3868 = ~n3854 & n3867;
  assign n3869 = ~n1481 & ~n3612;
  assign n3870 = n3261 & n3869;
  assign n3871 = n1466 & n3870;
  assign n3872 = x593 & n3580;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3605 & ~n3835;
  assign n3875 = x314 & x1050;
  assign n3876 = ~n3874 & n3875;
  assign n3877 = n2322 & n3346;
  assign n3878 = n3877 ^ x99;
  assign n3879 = n2634 & n3878;
  assign n3880 = x152 & n3372;
  assign n3881 = x161 & n3880;
  assign n3882 = x174 & n3370;
  assign n3883 = x144 & n3882;
  assign n3884 = ~n3881 & ~n3883;
  assign n3885 = n3353 & ~n3884;
  assign n3886 = ~n3879 & ~n3885;
  assign n3887 = n1496 & ~n2389;
  assign n3888 = x683 & ~n3887;
  assign n3889 = ~n2928 & ~n3888;
  assign n3890 = n2650 & n3889;
  assign n3891 = n2931 & ~n3890;
  assign n3892 = n2473 & ~n3891;
  assign n3893 = n1478 & n2935;
  assign n3894 = ~n2934 & n3893;
  assign n3895 = ~n3892 & ~n3894;
  assign n3896 = n2472 & ~n3895;
  assign n3897 = n3346 ^ x101;
  assign n3898 = n2634 & n3897;
  assign n3899 = ~x161 & n3880;
  assign n3900 = ~x144 & n3882;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = n3353 & ~n3901;
  assign n3903 = ~n3898 & ~n3902;
  assign n3904 = x65 & n3270;
  assign n3905 = n1752 & ~n2431;
  assign n3906 = ~n2865 & n3802;
  assign n3907 = ~x94 & x110;
  assign n3908 = n3459 & n3907;
  assign n3909 = ~n3242 & n3908;
  assign n3910 = ~n3906 & ~n3909;
  assign n3911 = x106 & n3442;
  assign n3912 = ~x24 & n3495;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = ~x999 & n3539;
  assign n3915 = ~n2565 & ~n3751;
  assign n3916 = x108 & ~n3282;
  assign n3917 = ~x98 & ~n3916;
  assign n3918 = n3448 & ~n3917;
  assign n3919 = ~n3915 & ~n3918;
  assign n3920 = n3448 & n3638;
  assign n3921 = n2426 & n3469;
  assign n3922 = x314 & n3921;
  assign n3923 = n3242 & n3908;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~x24 & n1572;
  assign n3926 = n3599 & n3925;
  assign n3927 = ~x314 & n3921;
  assign n3928 = ~n3926 & ~n3927;
  assign n3929 = x124 & ~x468;
  assign n3930 = n2323 & n3346;
  assign n3931 = n3930 ^ x113;
  assign n3932 = n2634 & n3931;
  assign n3933 = n3366 ^ x114;
  assign n3934 = n2634 & n3933;
  assign n3935 = ~x116 & n3365;
  assign n3936 = n3935 ^ x115;
  assign n3937 = n2634 & n3936;
  assign n3938 = n3365 ^ x116;
  assign n3939 = n2634 & n3938;
  assign n3940 = ~x87 & n2643;
  assign n3941 = n2973 & n3940;
  assign n3942 = x92 ^ x39;
  assign n3943 = x190 & n2481;
  assign n3944 = x178 & n2385;
  assign n3945 = ~n3943 & ~n3944;
  assign n3946 = n2980 & ~n3945;
  assign n3947 = x168 & n2481;
  assign n3948 = x157 & n2385;
  assign n3949 = ~n3947 & ~n3948;
  assign n3950 = n2982 & ~n3949;
  assign n3951 = ~n3946 & ~n3950;
  assign n3952 = n3951 ^ x92;
  assign n3953 = n3952 ^ n3951;
  assign n3954 = x178 ^ x157;
  assign n3955 = ~x299 & n3954;
  assign n3956 = n3955 ^ x157;
  assign n3957 = n3956 ^ n3951;
  assign n3958 = n3953 & ~n3957;
  assign n3959 = n3958 ^ n3951;
  assign n3960 = n3942 & ~n3959;
  assign n3961 = n3941 & n3960;
  assign n3962 = n2963 & ~n3961;
  assign n3963 = n1567 & ~n2952;
  assign n3987 = x173 ^ x151;
  assign n3988 = ~x299 & n3987;
  assign n3989 = n3988 ^ x151;
  assign n3990 = n3037 & ~n3989;
  assign n3991 = n2643 & ~n3990;
  assign n3992 = ~n2443 & ~n3991;
  assign n3993 = ~x150 & ~n3055;
  assign n3994 = x73 & ~x168;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = x299 & ~n3995;
  assign n3997 = ~x73 & x232;
  assign n3998 = n1205 & n3997;
  assign n3999 = n3055 & ~n3998;
  assign n4000 = ~x185 & ~x299;
  assign n4001 = ~n3999 & n4000;
  assign n4002 = x73 & ~x299;
  assign n4003 = ~x190 & n4002;
  assign n4004 = ~n4001 & ~n4003;
  assign n4005 = ~n3996 & n4004;
  assign n4006 = ~n3992 & n4005;
  assign n3964 = ~x54 & n1562;
  assign n3965 = ~n1565 & ~n1590;
  assign n3966 = n3964 & ~n3965;
  assign n3967 = x39 ^ x38;
  assign n3968 = n2975 ^ x38;
  assign n3969 = n2975 ^ x92;
  assign n3970 = ~n2975 & n3969;
  assign n3971 = n3970 ^ n2975;
  assign n3972 = n3968 & ~n3971;
  assign n3973 = n3972 ^ n3970;
  assign n3974 = n3973 ^ n2975;
  assign n3975 = n3974 ^ x92;
  assign n3976 = n3967 & n3975;
  assign n3977 = n3976 ^ x92;
  assign n3978 = n3966 & n3977;
  assign n3979 = n1574 & n3978;
  assign n3980 = ~x954 & n2958;
  assign n3981 = ~n2955 & n3980;
  assign n3982 = ~x79 & n3642;
  assign n3983 = x118 & ~n3982;
  assign n3984 = ~n3981 & ~n3983;
  assign n3985 = n1564 & ~n3984;
  assign n3986 = ~n3979 & ~n3985;
  assign n4007 = n4006 ^ n3986;
  assign n4008 = n3963 & n4007;
  assign n4009 = n4008 ^ n3986;
  assign n4010 = n3962 & ~n4009;
  assign n4011 = ~x163 & ~n3715;
  assign n4012 = n4011 ^ x150;
  assign n4013 = n3027 & ~n4012;
  assign n4014 = n1562 & ~n3078;
  assign n4015 = x165 & n2643;
  assign n4016 = n4014 & ~n4015;
  assign n4017 = ~n4013 & ~n4016;
  assign n4018 = ~n1729 & ~n4017;
  assign n4019 = ~n2643 & n4014;
  assign n4020 = n1569 & ~n4019;
  assign n4021 = ~n4018 & n4020;
  assign n4022 = ~x184 & ~n3719;
  assign n4023 = n4022 ^ x185;
  assign n4024 = n3027 & ~n4023;
  assign n4025 = ~x143 & n3725;
  assign n4026 = ~n4024 & ~n4025;
  assign n4027 = ~x299 & ~n4026;
  assign n4028 = n4021 & ~n4027;
  assign n4029 = ~n4010 & n4028;
  assign n4030 = x150 & n2643;
  assign n4031 = n4030 ^ n3984;
  assign n4032 = n3081 & n4031;
  assign n4033 = n4032 ^ n3984;
  assign n4034 = n3080 & ~n4033;
  assign n4035 = ~n1571 & n4017;
  assign n4036 = ~n4034 & n4035;
  assign n4037 = ~n4029 & ~n4036;
  assign n4038 = ~x109 & n1237;
  assign n4039 = n1303 & ~n4038;
  assign n4040 = ~n2469 & n4039;
  assign n4041 = n1305 & ~n1485;
  assign n4042 = ~n4040 & n4041;
  assign n4043 = n1752 & ~n4042;
  assign n4044 = n1678 & n2472;
  assign n4045 = ~n2666 & n3572;
  assign n4046 = ~n3835 & ~n4045;
  assign n4047 = ~n4044 & n4046;
  assign n4048 = ~n4043 & n4047;
  assign n4049 = n4048 ^ x128;
  assign n4050 = ~x228 & ~n4049;
  assign n4051 = n4050 ^ x128;
  assign n4052 = n1571 & ~n2681;
  assign n4053 = ~n2642 & n4052;
  assign n4054 = ~n2901 & ~n4053;
  assign n4055 = ~x31 & ~x80;
  assign n4056 = x818 & n4055;
  assign n4057 = x1093 & n4056;
  assign n4058 = x951 & x982;
  assign n4059 = n2868 & n4058;
  assign n4060 = n2872 & n4059;
  assign n4061 = ~n4057 & ~n4060;
  assign n4062 = ~x120 & n4061;
  assign n4063 = n4054 & ~n4062;
  assign n4064 = ~x24 & n3638;
  assign n4065 = n3044 & n4064;
  assign n4066 = n2435 & n4065;
  assign n4067 = x181 & n2364;
  assign n4068 = x159 & n2367;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = n3292 & ~n4069;
  assign n4071 = ~n3354 & ~n3357;
  assign n4072 = n2565 & ~n4071;
  assign n4073 = ~n2566 & ~n4072;
  assign n4074 = ~x146 & ~n1729;
  assign n4075 = n1490 & n1571;
  assign n4076 = x51 & ~x87;
  assign n4077 = ~n4075 & n4076;
  assign n4078 = ~n4074 & n4077;
  assign n4079 = n1729 ^ x163;
  assign n4080 = n4079 ^ x163;
  assign n4081 = x184 ^ x163;
  assign n4082 = n4080 & n4081;
  assign n4083 = n4082 ^ x163;
  assign n4084 = x87 & ~n4083;
  assign n4085 = ~n4078 & ~n4084;
  assign n4086 = n4073 & n4085;
  assign n4087 = ~n4070 & ~n4086;
  assign n4088 = ~n4066 & n4087;
  assign n4089 = n2643 & ~n4088;
  assign n4097 = n3703 & ~n4064;
  assign n4090 = x24 & x77;
  assign n4091 = ~x86 & ~n4090;
  assign n4092 = ~n3638 & n4091;
  assign n4093 = ~x39 & ~n4092;
  assign n4094 = n2561 & n4093;
  assign n4095 = n1468 & n4094;
  assign n4096 = n1444 & n4095;
  assign n4098 = n4097 ^ n4096;
  assign n4099 = n4098 ^ n4097;
  assign n4100 = x72 ^ x39;
  assign n4101 = n2562 & n4100;
  assign n4102 = x39 & n2482;
  assign n4103 = n4101 & ~n4102;
  assign n4104 = ~x125 & ~x133;
  assign n4105 = n4104 ^ x121;
  assign n4106 = ~x134 & ~x135;
  assign n4107 = ~x136 & n4106;
  assign n4108 = ~x130 & n4107;
  assign n4109 = ~x126 & ~x132;
  assign n4110 = n4108 & n4109;
  assign n4111 = n4104 & n4110;
  assign n4112 = n4105 & n4111;
  assign n4113 = n4112 ^ n4105;
  assign n4114 = ~n4103 & ~n4113;
  assign n4115 = n4114 ^ n4097;
  assign n4116 = ~n4099 & n4115;
  assign n4117 = n4116 ^ n4097;
  assign n4118 = n2566 & n4117;
  assign n4119 = ~n4089 & ~n4118;
  assign n4120 = ~x90 & ~x111;
  assign n4121 = ~x72 & n4120;
  assign n4122 = n2424 & n4121;
  assign n4123 = n2435 & ~n4122;
  assign n4124 = x39 & ~x110;
  assign n4125 = n2573 & n4124;
  assign n4126 = n2643 & ~n3417;
  assign n4127 = ~x39 & x110;
  assign n4128 = n2389 & n4127;
  assign n4129 = ~n2331 & n4128;
  assign n4130 = ~n4126 & n4129;
  assign n4131 = ~n4125 & ~n4130;
  assign n4132 = ~n4123 & n4131;
  assign n4133 = ~n1455 & ~n4092;
  assign n4134 = ~x39 & ~n3599;
  assign n4135 = ~n4133 & n4134;
  assign n4136 = n2560 & ~n4135;
  assign n4137 = ~x287 & n2643;
  assign n4138 = x158 & n1737;
  assign n4139 = n4137 & n4138;
  assign n4140 = n2669 & ~n4139;
  assign n4141 = n1574 & ~n4140;
  assign n4142 = n1232 ^ x172;
  assign n4143 = n4142 ^ x172;
  assign n4144 = x172 ^ x152;
  assign n4145 = n4144 ^ x172;
  assign n4146 = ~n4143 & ~n4145;
  assign n4147 = n4146 ^ x172;
  assign n4148 = ~x51 & n4147;
  assign n4149 = n4148 ^ x172;
  assign n4150 = x299 & ~n4149;
  assign n4151 = n2643 & ~n4150;
  assign n4152 = ~n4141 & ~n4151;
  assign n4153 = ~x72 & n2559;
  assign n4154 = x180 & ~x287;
  assign n4155 = n2346 & n4154;
  assign n4156 = x224 & ~n4155;
  assign n4157 = ~x51 & x222;
  assign n4158 = ~x223 & n4157;
  assign n4159 = n1232 & n4158;
  assign n4160 = ~n4156 & n4159;
  assign n4161 = n4153 & n4160;
  assign n4162 = x193 ^ x51;
  assign n4163 = n4162 ^ x193;
  assign n4164 = n4163 ^ x299;
  assign n4165 = n1232 ^ x174;
  assign n4166 = ~x174 & n4165;
  assign n4167 = n4166 ^ x193;
  assign n4168 = n4167 ^ x174;
  assign n4169 = n4164 & ~n4168;
  assign n4170 = n4169 ^ n4166;
  assign n4171 = n4170 ^ x174;
  assign n4172 = ~x299 & ~n4171;
  assign n4173 = n4172 ^ x299;
  assign n4174 = ~n4161 & ~n4173;
  assign n4175 = ~n4152 & ~n4174;
  assign n4176 = x39 & ~n4175;
  assign n4177 = n4136 & ~n4176;
  assign n4178 = n4151 & n4173;
  assign n4179 = ~x121 & ~x125;
  assign n4180 = n4110 & n4179;
  assign n4181 = x133 ^ x125;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = n2566 & ~n4182;
  assign n4184 = ~n4178 & ~n4183;
  assign n4185 = ~n4177 & n4184;
  assign n4186 = x39 & n2560;
  assign n4187 = ~n2484 & n4186;
  assign n4188 = n4153 & n4187;
  assign n4189 = ~n4175 & n4188;
  assign n4190 = ~x87 & ~n4189;
  assign n4191 = ~n4185 & n4190;
  assign n4192 = x87 & n2643;
  assign n4193 = x162 ^ x140;
  assign n4194 = x299 & n4193;
  assign n4195 = n4194 ^ x140;
  assign n4196 = n4192 & n4195;
  assign n4197 = n1571 & ~n4196;
  assign n4198 = ~n4191 & n4197;
  assign n4199 = n1567 & n4096;
  assign n4200 = x197 ^ x145;
  assign n4201 = x299 & n4200;
  assign n4202 = n4201 ^ x145;
  assign n4203 = n4202 ^ n3135;
  assign n4204 = n4091 & n4203;
  assign n4205 = n4204 ^ n3135;
  assign n4206 = n2643 & n4205;
  assign n4207 = n4199 & ~n4206;
  assign n4208 = n3940 & n4149;
  assign n4209 = x162 & n4192;
  assign n4210 = ~n1571 & ~n4209;
  assign n4211 = ~n4208 & n4210;
  assign n4212 = ~n4183 & n4211;
  assign n4213 = ~n4207 & ~n4212;
  assign n4214 = ~n4198 & n4213;
  assign n4215 = ~x121 & n4104;
  assign n4216 = n4215 ^ x126;
  assign n4217 = n2566 & n4216;
  assign n4218 = ~n4110 & n4217;
  assign n4219 = ~n4199 & ~n4218;
  assign n4220 = ~n4103 & ~n4219;
  assign n4221 = x160 & n4137;
  assign n4222 = n2367 & ~n4221;
  assign n4223 = x182 & n4137;
  assign n4224 = n2364 & ~n4223;
  assign n4225 = ~n4222 & ~n4224;
  assign n4226 = n2564 & ~n4225;
  assign n4227 = x166 ^ x153;
  assign n4228 = ~x51 & ~n4227;
  assign n4229 = n4228 ^ x153;
  assign n4230 = n3940 & n4229;
  assign n4231 = ~n1571 & n4230;
  assign n4232 = ~n2566 & ~n4231;
  assign n4233 = ~n4226 & ~n4232;
  assign n4234 = ~n4220 & n4233;
  assign n4235 = n3956 ^ n3151;
  assign n4236 = ~n4091 & n4235;
  assign n4237 = n4236 ^ n3151;
  assign n4238 = n4199 & n4237;
  assign n4241 = x185 ^ x150;
  assign n4239 = x299 ^ x150;
  assign n4240 = n4239 ^ x150;
  assign n4242 = n4241 ^ n4240;
  assign n4243 = n1571 ^ x150;
  assign n4244 = n4243 ^ x150;
  assign n4245 = n4244 ^ n4240;
  assign n4246 = ~n4240 & ~n4245;
  assign n4247 = n4246 ^ n4240;
  assign n4248 = ~n4242 & ~n4247;
  assign n4249 = n4248 ^ n4246;
  assign n4250 = n4249 ^ x150;
  assign n4251 = n4250 ^ n4240;
  assign n4252 = n4251 ^ n1571;
  assign n4253 = n4252 ^ n4251;
  assign n4254 = x299 ^ x153;
  assign n4255 = n4254 ^ x153;
  assign n4256 = x175 ^ x153;
  assign n4257 = ~n4255 & n4256;
  assign n4258 = n4257 ^ x153;
  assign n4259 = n4258 ^ n1232;
  assign n4260 = n4259 ^ n4258;
  assign n4261 = n4258 ^ n3665;
  assign n4262 = n4261 ^ n4258;
  assign n4263 = ~n4260 & ~n4262;
  assign n4264 = n4263 ^ n4258;
  assign n4265 = ~x51 & n4264;
  assign n4266 = n4265 ^ n4258;
  assign n4267 = n4266 ^ n4251;
  assign n4268 = n4267 ^ n4251;
  assign n4269 = n4253 & n4268;
  assign n4270 = n4269 ^ n4251;
  assign n4271 = ~x87 & ~n4270;
  assign n4272 = n4271 ^ n4251;
  assign n4273 = ~n4238 & n4272;
  assign n4274 = n2643 & ~n4273;
  assign n4275 = ~n4234 & ~n4274;
  assign n4276 = x250 & n2651;
  assign n4277 = n4276 ^ x127;
  assign n4278 = n4277 ^ x127;
  assign n4279 = n2320 ^ x127;
  assign n4280 = n4278 & n4279;
  assign n4281 = n4280 ^ x127;
  assign n4282 = x94 & ~n4281;
  assign n4283 = x129 & ~n4282;
  assign n4284 = ~n3751 & n4283;
  assign n4285 = ~x100 & ~n2651;
  assign n4286 = ~x250 & ~n4285;
  assign n4287 = n4286 ^ x129;
  assign n4288 = n4287 ^ x129;
  assign n4289 = n2929 & n4288;
  assign n4290 = n4289 ^ x129;
  assign n4291 = ~n1561 & ~n4290;
  assign n4292 = ~n1632 & ~n4291;
  assign n4293 = ~n1752 & ~n4292;
  assign n4294 = x140 & n1775;
  assign n4295 = n1737 & n3147;
  assign n4296 = ~n4294 & ~n4295;
  assign n4297 = n4137 & ~n4296;
  assign n4298 = n2669 & ~n4297;
  assign n4299 = n1574 & ~n4298;
  assign n4300 = x39 & ~n4299;
  assign n4301 = n4136 & ~n4300;
  assign n4302 = ~x87 & n1571;
  assign n4303 = n4109 & n4215;
  assign n4304 = n4303 ^ x130;
  assign n4305 = n4303 ^ n4107;
  assign n4306 = n4303 ^ n1232;
  assign n4307 = n4303 & n4306;
  assign n4308 = n4307 ^ n4303;
  assign n4309 = n4305 & n4308;
  assign n4310 = n4309 ^ n4307;
  assign n4311 = n4310 ^ n4303;
  assign n4312 = n4311 ^ n1232;
  assign n4313 = n4304 & n4312;
  assign n4314 = n4313 ^ n1232;
  assign n4315 = ~n4188 & n4314;
  assign n4316 = ~n1232 & n3023;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = n4302 & n4317;
  assign n4319 = ~n4301 & n4318;
  assign n4320 = ~n1232 & n2643;
  assign n4321 = x169 & n4320;
  assign n4322 = ~n1571 & ~n4192;
  assign n4323 = ~n4321 & n4322;
  assign n4324 = ~n4314 & n4323;
  assign n4325 = ~n4319 & ~n4324;
  assign n4326 = ~x51 & ~n4325;
  assign n4327 = n1729 ^ x188;
  assign n4328 = n4327 ^ x188;
  assign n4329 = n3164 & ~n4328;
  assign n4330 = n4329 ^ x188;
  assign n4331 = n2643 & n4330;
  assign n4332 = x87 & ~n4331;
  assign n4333 = ~n4326 & ~n4332;
  assign n4334 = ~n2484 & n2564;
  assign n4335 = n2566 & ~n4334;
  assign n4336 = ~n4096 & n4335;
  assign n4337 = n2643 & n3670;
  assign n4338 = ~x24 & x77;
  assign n4339 = ~n4337 & n4338;
  assign n4340 = x149 & n2366;
  assign n4341 = x183 & n1775;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~n4339 & ~n4342;
  assign n4344 = n4137 & n4343;
  assign n4345 = n2566 & n4344;
  assign n4346 = ~n4336 & ~n4345;
  assign n4347 = n4108 ^ x132;
  assign n4348 = x132 ^ x126;
  assign n4349 = ~x132 & n4348;
  assign n4350 = n4349 ^ x132;
  assign n4351 = ~n4347 & ~n4350;
  assign n4352 = n4351 ^ n4349;
  assign n4353 = n4352 ^ x132;
  assign n4354 = n4353 ^ x126;
  assign n4355 = n4215 & n4354;
  assign n4356 = n4355 ^ x132;
  assign n4357 = ~n4103 & n4356;
  assign n4358 = ~n4346 & ~n4357;
  assign n4359 = n4199 & ~n4339;
  assign n4360 = n1729 ^ x190;
  assign n4361 = n4360 ^ x190;
  assign n4362 = x190 ^ x168;
  assign n4363 = ~n4361 & n4362;
  assign n4364 = n4363 ^ x190;
  assign n4365 = ~n1232 & n4364;
  assign n4366 = n2565 & ~n4365;
  assign n4367 = x299 ^ x164;
  assign n4368 = n4367 ^ x164;
  assign n4369 = n4368 ^ n2965;
  assign n4370 = n1571 ^ x164;
  assign n4371 = n4370 ^ x164;
  assign n4372 = n4371 ^ n4368;
  assign n4373 = ~n4368 & ~n4372;
  assign n4374 = n4373 ^ n4368;
  assign n4375 = ~n4369 & ~n4374;
  assign n4376 = n4375 ^ n4373;
  assign n4377 = n4376 ^ x164;
  assign n4378 = n4377 ^ n4368;
  assign n4379 = x87 & n4378;
  assign n4380 = n2643 & ~n4379;
  assign n4381 = n1729 ^ x173;
  assign n4382 = n4381 ^ x173;
  assign n4383 = n3987 & ~n4382;
  assign n4384 = n4383 ^ x173;
  assign n4385 = n4076 & ~n4384;
  assign n4386 = n4380 & ~n4385;
  assign n4387 = ~n4366 & n4386;
  assign n4388 = ~n4359 & ~n4387;
  assign n4389 = ~n4358 & n4388;
  assign n4390 = x145 & n1775;
  assign n4391 = x197 & n2366;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = n4137 & ~n4392;
  assign n4394 = ~x72 & n2669;
  assign n4395 = ~n4393 & n4394;
  assign n4396 = n4100 & ~n4395;
  assign n4397 = ~n3751 & n4396;
  assign n4400 = ~x133 & ~n4180;
  assign n4401 = n4335 & ~n4400;
  assign n4402 = n1729 ^ x183;
  assign n4403 = n4402 ^ x183;
  assign n4404 = x183 ^ x149;
  assign n4405 = ~n4403 & n4404;
  assign n4406 = n4405 ^ x183;
  assign n4407 = n4192 & n4406;
  assign n4408 = ~n4401 & ~n4407;
  assign n4398 = ~x86 & n2918;
  assign n4399 = ~n3004 & ~n4398;
  assign n4409 = n4408 ^ n4399;
  assign n4410 = ~n4199 & n4409;
  assign n4411 = n4410 ^ n4399;
  assign n4412 = ~n4397 & n4411;
  assign n4413 = n2565 & ~n4096;
  assign n4426 = x192 ^ x171;
  assign n4427 = n1729 & n4426;
  assign n4428 = n4427 ^ x171;
  assign n4414 = ~x130 & n4303;
  assign n4415 = ~x136 & n4414;
  assign n4416 = ~x135 & n4415;
  assign n4417 = x134 & ~n4416;
  assign n4418 = ~n4103 & ~n4417;
  assign n4419 = x186 & n1775;
  assign n4420 = x164 & n2366;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = n4137 & ~n4421;
  assign n4423 = n4394 & ~n4422;
  assign n4424 = n4101 & ~n4423;
  assign n4425 = ~n4418 & ~n4424;
  assign n4429 = n4428 ^ n4425;
  assign n4430 = n4429 ^ n4425;
  assign n4431 = n4425 ^ n2643;
  assign n4432 = n4431 ^ n4425;
  assign n4433 = n4430 & n4432;
  assign n4434 = n4433 ^ n4425;
  assign n4435 = ~n1232 & ~n4434;
  assign n4436 = n4435 ^ n4425;
  assign n4437 = n4413 & n4436;
  assign n4438 = x150 & n2366;
  assign n4439 = x185 & n1775;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = n4137 & ~n4440;
  assign n4442 = n4334 & ~n4441;
  assign n4443 = n1232 & ~n4442;
  assign n4445 = ~x134 & n4416;
  assign n4444 = n4415 ^ x135;
  assign n4446 = n4445 ^ n4444;
  assign n4447 = ~n4103 & n4446;
  assign n4448 = n4443 & ~n4447;
  assign n4449 = x194 ^ x170;
  assign n4450 = n1729 & n4449;
  assign n4451 = n4450 ^ x170;
  assign n4452 = n4320 & n4451;
  assign n4453 = ~n4448 & ~n4452;
  assign n4454 = n4413 & n4453;
  assign n4455 = x163 & n2366;
  assign n4456 = x184 & n1775;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = n4137 & ~n4457;
  assign n4459 = n2669 & ~n4458;
  assign n4460 = n4153 & ~n4459;
  assign n4461 = x39 & n1232;
  assign n4462 = ~n4460 & n4461;
  assign n4463 = n2643 & n3171;
  assign n4464 = ~n1232 & ~n4463;
  assign n4465 = n2561 & ~n4464;
  assign n4466 = ~n4462 & n4465;
  assign n4467 = ~n4135 & n4466;
  assign n4473 = n4414 ^ x136;
  assign n4468 = n1729 ^ x148;
  assign n4469 = n4468 ^ x148;
  assign n4470 = n3169 & n4469;
  assign n4471 = n4470 ^ x148;
  assign n4472 = n4320 & n4471;
  assign n4474 = n4473 ^ n4472;
  assign n4475 = n4472 ^ n1232;
  assign n4476 = n4475 ^ n4472;
  assign n4477 = n4474 & n4476;
  assign n4478 = ~n4107 & n4477;
  assign n4479 = n4478 ^ n4475;
  assign n4480 = ~n4334 & n4479;
  assign n4481 = n2565 & ~n4480;
  assign n4482 = ~n4467 & n4481;
  assign n4483 = ~x198 & n3415;
  assign n4484 = ~x210 & n3416;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = n2978 & ~n4485;
  assign n4487 = ~n3377 & n4486;
  assign n4488 = ~x39 & x137;
  assign n4489 = ~n4487 & ~n4488;
  assign n4490 = n2953 ^ x138;
  assign n4491 = x139 ^ x138;
  assign n4492 = ~x138 & n4491;
  assign n4493 = n4492 ^ x138;
  assign n4494 = ~n4490 & ~n4493;
  assign n4495 = n4494 ^ n4492;
  assign n4496 = n4495 ^ x138;
  assign n4497 = n4496 ^ x139;
  assign n4498 = n3980 & n4497;
  assign n4499 = n4498 ^ x138;
  assign n4500 = n4499 ^ n4463;
  assign n4501 = n4500 ^ n4463;
  assign n4502 = n1565 & n1569;
  assign n4503 = n2973 ^ n2948;
  assign n4504 = n4503 ^ n2948;
  assign n4505 = n2948 ^ n2386;
  assign n4506 = n4505 ^ n2948;
  assign n4507 = n4504 & n4506;
  assign n4508 = n4507 ^ n2948;
  assign n4509 = x39 & ~n4508;
  assign n4510 = n4509 ^ n2948;
  assign n4511 = n4502 & ~n4510;
  assign n4512 = n1615 & n3080;
  assign n4513 = ~n4511 & n4512;
  assign n4514 = n4513 ^ n4463;
  assign n4515 = n4514 ^ n4463;
  assign n4516 = n4501 & n4515;
  assign n4517 = n4516 ^ n4463;
  assign n4518 = n3607 & ~n4517;
  assign n4519 = n4518 ^ n4463;
  assign n4520 = n3980 ^ x139;
  assign n4521 = ~n2955 & n4520;
  assign n4522 = n4521 ^ n3023;
  assign n4523 = n4522 ^ n3023;
  assign n4524 = n4513 ^ n3023;
  assign n4525 = n4524 ^ n3023;
  assign n4526 = n4523 & n4525;
  assign n4527 = n4526 ^ n3023;
  assign n4528 = n3607 & ~n4527;
  assign n4529 = n4528 ^ n3023;
  assign n4530 = ~n2390 & n3290;
  assign n4531 = x35 & ~x93;
  assign n4532 = ~x841 & n4531;
  assign n4533 = n1450 & n4532;
  assign n4534 = ~x45 & ~x47;
  assign n4535 = ~x102 & n4534;
  assign n4536 = ~n3281 & n4535;
  assign n4537 = ~n4533 & n4536;
  assign n4538 = ~x47 & ~n1229;
  assign n4539 = ~x252 & ~n4538;
  assign n4540 = ~n4537 & ~n4539;
  assign n4541 = ~x40 & ~n4540;
  assign n4542 = ~n4530 & n4541;
  assign n4543 = n3598 & n4542;
  assign n4544 = ~n3751 & ~n4543;
  assign n4545 = ~n2666 & ~n3573;
  assign n4546 = ~x287 & ~n3295;
  assign n4547 = ~x120 & ~n4546;
  assign n4548 = ~n2397 & ~n4547;
  assign n4549 = n2567 & n4548;
  assign n4550 = ~n4545 & ~n4549;
  assign n4551 = ~n4544 & n4550;
  assign n4552 = n2868 & ~n4551;
  assign n4553 = x832 & n2868;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = x1154 ^ x618;
  assign n4556 = x781 & n4555;
  assign n4557 = x1155 ^ x609;
  assign n4558 = x785 & n4557;
  assign n4559 = ~n4556 & ~n4558;
  assign n4560 = x1157 ^ x630;
  assign n4561 = x787 & n4560;
  assign n4562 = x1158 ^ x626;
  assign n4563 = x788 & n4562;
  assign n4564 = ~n4561 & ~n4563;
  assign n4565 = n4559 & n4564;
  assign n4566 = x1160 ^ x644;
  assign n4567 = x790 & n4566;
  assign n4568 = x603 & ~n4567;
  assign n4569 = n4565 & n4568;
  assign n4570 = x1159 ^ x619;
  assign n4571 = x789 & n4570;
  assign n4572 = x1153 ^ x608;
  assign n4573 = x778 & n4572;
  assign n4574 = ~n4571 & ~n4573;
  assign n4575 = x1156 ^ x629;
  assign n4576 = x792 & n4575;
  assign n4577 = n4574 & ~n4576;
  assign n4578 = n4569 & n4577;
  assign n4579 = x621 & x1091;
  assign n4580 = n4578 & ~n4579;
  assign n4581 = x1160 ^ x715;
  assign n4582 = x790 & n4581;
  assign n4583 = x1158 ^ x641;
  assign n4584 = x788 & n4583;
  assign n4585 = ~n4582 & ~n4584;
  assign n4586 = x1153 ^ x625;
  assign n4587 = x778 & n4586;
  assign n4588 = n4585 & ~n4587;
  assign n4589 = x1155 ^ x660;
  assign n4590 = x785 & n4589;
  assign n4591 = x680 & ~n4590;
  assign n4592 = x1154 ^ x627;
  assign n4593 = x781 & n4592;
  assign n4594 = x1157 ^ x647;
  assign n4595 = x787 & n4594;
  assign n4596 = ~n4593 & ~n4595;
  assign n4597 = n4591 & n4596;
  assign n4598 = n4588 & n4597;
  assign n4599 = x1156 ^ x628;
  assign n4600 = x792 & n4599;
  assign n4601 = x1159 ^ x648;
  assign n4602 = x789 & n4601;
  assign n4603 = ~n4600 & ~n4602;
  assign n4604 = n4598 & n4603;
  assign n4605 = x665 & x1091;
  assign n4606 = n4604 & ~n4605;
  assign n4607 = n4606 ^ x761;
  assign n4608 = n4607 ^ x761;
  assign n4609 = x761 ^ x738;
  assign n4610 = n4609 ^ x761;
  assign n4611 = n4608 & ~n4610;
  assign n4612 = n4611 ^ x761;
  assign n4613 = ~n4580 & ~n4612;
  assign n4614 = n4613 ^ x761;
  assign n4615 = n4614 ^ x140;
  assign n4616 = ~n4554 & n4615;
  assign n4617 = n4616 ^ x140;
  assign n4618 = n4606 ^ x749;
  assign n4619 = n4618 ^ x749;
  assign n4620 = x749 ^ x706;
  assign n4621 = n4620 ^ x749;
  assign n4622 = n4619 & n4621;
  assign n4623 = n4622 ^ x749;
  assign n4624 = ~n4580 & n4623;
  assign n4625 = n4624 ^ x749;
  assign n4626 = n4625 ^ x141;
  assign n4627 = ~n4554 & ~n4626;
  assign n4628 = n4627 ^ x141;
  assign n4629 = x743 ^ x735;
  assign n4630 = n4629 ^ x743;
  assign n4631 = n4606 ^ x743;
  assign n4632 = n4631 ^ x743;
  assign n4633 = n4630 & n4632;
  assign n4634 = n4633 ^ x743;
  assign n4635 = ~n4580 & n4634;
  assign n4636 = n4635 ^ x743;
  assign n4637 = n4636 ^ x142;
  assign n4638 = ~n4554 & n4637;
  assign n4639 = n4638 ^ x142;
  assign n4640 = n4606 ^ x774;
  assign n4641 = n4640 ^ x774;
  assign n4642 = x774 ^ x687;
  assign n4643 = n4642 ^ x774;
  assign n4644 = n4641 & n4643;
  assign n4645 = n4644 ^ x774;
  assign n4646 = ~n4580 & ~n4645;
  assign n4647 = n4646 ^ x774;
  assign n4648 = n4647 ^ x143;
  assign n4649 = ~n4554 & n4648;
  assign n4650 = n4649 ^ x143;
  assign n4651 = n4606 ^ x758;
  assign n4652 = n4651 ^ x758;
  assign n4653 = x758 ^ x736;
  assign n4654 = n4653 ^ x758;
  assign n4655 = n4652 & n4654;
  assign n4656 = n4655 ^ x758;
  assign n4657 = ~n4580 & n4656;
  assign n4658 = n4657 ^ x758;
  assign n4659 = n4658 ^ x144;
  assign n4660 = ~n4554 & n4659;
  assign n4661 = n4660 ^ x144;
  assign n4662 = n4606 ^ x767;
  assign n4663 = n4662 ^ x767;
  assign n4664 = x767 ^ x698;
  assign n4665 = n4664 ^ x767;
  assign n4666 = n4663 & ~n4665;
  assign n4667 = n4666 ^ x767;
  assign n4668 = ~n4580 & ~n4667;
  assign n4669 = n4668 ^ x767;
  assign n4670 = n4669 ^ x145;
  assign n4671 = ~n4554 & n4670;
  assign n4672 = n4671 ^ x145;
  assign n4673 = x907 ^ x743;
  assign n4674 = n4673 ^ x743;
  assign n4675 = n4630 & n4674;
  assign n4676 = n4675 ^ x743;
  assign n4677 = ~x947 & n4676;
  assign n4678 = n4677 ^ x743;
  assign n4679 = n4678 ^ x146;
  assign n4680 = ~n4554 & n4679;
  assign n4681 = n4680 ^ x146;
  assign n4682 = x770 ^ x726;
  assign n4683 = n4682 ^ x770;
  assign n4684 = x907 ^ x770;
  assign n4685 = n4684 ^ x770;
  assign n4686 = n4683 & n4685;
  assign n4687 = n4686 ^ x770;
  assign n4688 = ~x947 & ~n4687;
  assign n4689 = n4688 ^ x770;
  assign n4690 = n4689 ^ x147;
  assign n4691 = ~n4554 & n4690;
  assign n4692 = n4691 ^ x147;
  assign n4693 = x907 ^ x749;
  assign n4694 = n4693 ^ x749;
  assign n4695 = n4621 & n4694;
  assign n4696 = n4695 ^ x749;
  assign n4697 = ~x947 & n4696;
  assign n4698 = n4697 ^ x749;
  assign n4699 = n4698 ^ x148;
  assign n4700 = ~n4554 & ~n4699;
  assign n4701 = n4700 ^ x148;
  assign n4702 = ~n2394 & ~n4547;
  assign n4703 = n2392 & n2664;
  assign n4704 = n2663 & ~n2974;
  assign n4705 = ~n4703 & ~n4704;
  assign n4706 = ~n4702 & n4705;
  assign n4707 = n2567 & ~n4706;
  assign n4708 = ~n4544 & ~n4707;
  assign n4709 = n2868 & ~n4708;
  assign n4710 = ~n4553 & ~n4709;
  assign n4711 = x755 ^ x725;
  assign n4712 = n4711 ^ x755;
  assign n4713 = x907 ^ x755;
  assign n4714 = n4713 ^ x755;
  assign n4715 = ~n4712 & n4714;
  assign n4716 = n4715 ^ x755;
  assign n4717 = ~x947 & ~n4716;
  assign n4718 = n4717 ^ x755;
  assign n4719 = ~n4710 & ~n4718;
  assign n4720 = ~x149 & n4554;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = x751 ^ x701;
  assign n4723 = n4722 ^ x751;
  assign n4724 = x907 ^ x751;
  assign n4725 = n4724 ^ x751;
  assign n4726 = ~n4723 & n4725;
  assign n4727 = n4726 ^ x751;
  assign n4728 = ~x947 & ~n4727;
  assign n4729 = n4728 ^ x751;
  assign n4730 = ~n4710 & ~n4729;
  assign n4731 = ~x150 & n4554;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733 = x745 ^ x723;
  assign n4734 = n4733 ^ x745;
  assign n4735 = x907 ^ x745;
  assign n4736 = n4735 ^ x745;
  assign n4737 = ~n4734 & n4736;
  assign n4738 = n4737 ^ x745;
  assign n4739 = ~x947 & ~n4738;
  assign n4740 = n4739 ^ x745;
  assign n4741 = n4740 ^ x151;
  assign n4742 = ~n4554 & n4741;
  assign n4743 = n4742 ^ x151;
  assign n4744 = x759 ^ x696;
  assign n4745 = n4744 ^ x759;
  assign n4746 = x907 ^ x759;
  assign n4747 = n4746 ^ x759;
  assign n4748 = n4745 & n4747;
  assign n4749 = n4748 ^ x759;
  assign n4750 = ~x947 & n4749;
  assign n4751 = n4750 ^ x759;
  assign n4752 = n4751 ^ x152;
  assign n4753 = ~n4554 & n4752;
  assign n4754 = n4753 ^ x152;
  assign n4755 = x766 ^ x700;
  assign n4756 = n4755 ^ x766;
  assign n4757 = x907 ^ x766;
  assign n4758 = n4757 ^ x766;
  assign n4759 = n4756 & n4758;
  assign n4760 = n4759 ^ x766;
  assign n4761 = ~x947 & n4760;
  assign n4762 = n4761 ^ x766;
  assign n4763 = n4762 ^ x153;
  assign n4764 = ~n4554 & ~n4763;
  assign n4765 = n4764 ^ x153;
  assign n4766 = x742 ^ x704;
  assign n4767 = n4766 ^ x742;
  assign n4768 = x907 ^ x742;
  assign n4769 = n4768 ^ x742;
  assign n4770 = ~n4767 & n4769;
  assign n4771 = n4770 ^ x742;
  assign n4772 = ~x947 & ~n4771;
  assign n4773 = n4772 ^ x742;
  assign n4774 = ~n4710 & ~n4773;
  assign n4775 = ~x154 & n4554;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = x757 ^ x686;
  assign n4778 = n4777 ^ x757;
  assign n4779 = x907 ^ x757;
  assign n4780 = n4779 ^ x757;
  assign n4781 = ~n4778 & n4780;
  assign n4782 = n4781 ^ x757;
  assign n4783 = ~x947 & ~n4782;
  assign n4784 = n4783 ^ x757;
  assign n4785 = ~n4710 & ~n4784;
  assign n4786 = ~x155 & n4554;
  assign n4787 = ~n4785 & ~n4786;
  assign n4788 = x741 ^ x724;
  assign n4789 = n4788 ^ x741;
  assign n4790 = x907 ^ x741;
  assign n4791 = n4790 ^ x741;
  assign n4792 = ~n4789 & n4791;
  assign n4793 = n4792 ^ x741;
  assign n4794 = ~x947 & ~n4793;
  assign n4795 = n4794 ^ x741;
  assign n4796 = ~n4710 & ~n4795;
  assign n4797 = ~x156 & n4554;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = x760 ^ x688;
  assign n4800 = n4799 ^ x760;
  assign n4801 = x907 ^ x760;
  assign n4802 = n4801 ^ x760;
  assign n4803 = ~n4800 & n4802;
  assign n4804 = n4803 ^ x760;
  assign n4805 = ~x947 & ~n4804;
  assign n4806 = n4805 ^ x760;
  assign n4807 = n4806 ^ x157;
  assign n4808 = ~n4554 & n4807;
  assign n4809 = n4808 ^ x157;
  assign n4810 = x753 ^ x702;
  assign n4811 = n4810 ^ x753;
  assign n4812 = x907 ^ x753;
  assign n4813 = n4812 ^ x753;
  assign n4814 = ~n4811 & n4813;
  assign n4815 = n4814 ^ x753;
  assign n4816 = ~x947 & ~n4815;
  assign n4817 = n4816 ^ x753;
  assign n4818 = ~n4710 & ~n4817;
  assign n4819 = ~x158 & n4554;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = x754 ^ x709;
  assign n4822 = n4821 ^ x754;
  assign n4823 = x907 ^ x754;
  assign n4824 = n4823 ^ x754;
  assign n4825 = ~n4822 & n4824;
  assign n4826 = n4825 ^ x754;
  assign n4827 = ~x947 & ~n4826;
  assign n4828 = n4827 ^ x754;
  assign n4829 = n4828 ^ x159;
  assign n4830 = ~n4554 & n4829;
  assign n4831 = n4830 ^ x159;
  assign n4832 = x756 ^ x734;
  assign n4833 = n4832 ^ x756;
  assign n4834 = x907 ^ x756;
  assign n4835 = n4834 ^ x756;
  assign n4836 = ~n4833 & n4835;
  assign n4837 = n4836 ^ x756;
  assign n4838 = ~x947 & ~n4837;
  assign n4839 = n4838 ^ x756;
  assign n4840 = n4839 ^ x160;
  assign n4841 = ~n4554 & n4840;
  assign n4842 = n4841 ^ x160;
  assign n4843 = x907 ^ x758;
  assign n4844 = n4843 ^ x758;
  assign n4845 = n4654 & n4844;
  assign n4846 = n4845 ^ x758;
  assign n4847 = ~x947 & n4846;
  assign n4848 = n4847 ^ x758;
  assign n4849 = n4848 ^ x161;
  assign n4850 = ~n4554 & n4849;
  assign n4851 = n4850 ^ x161;
  assign n4852 = x907 ^ x761;
  assign n4853 = n4852 ^ x761;
  assign n4854 = ~n4610 & n4853;
  assign n4855 = n4854 ^ x761;
  assign n4856 = ~x947 & ~n4855;
  assign n4857 = n4856 ^ x761;
  assign n4858 = n4857 ^ x162;
  assign n4859 = ~n4554 & n4858;
  assign n4860 = n4859 ^ x162;
  assign n4861 = x777 ^ x737;
  assign n4862 = n4861 ^ x777;
  assign n4863 = x907 ^ x777;
  assign n4864 = n4863 ^ x777;
  assign n4865 = ~n4862 & n4864;
  assign n4866 = n4865 ^ x777;
  assign n4867 = ~x947 & ~n4866;
  assign n4868 = n4867 ^ x777;
  assign n4869 = n4868 ^ x163;
  assign n4870 = ~n4554 & n4869;
  assign n4871 = n4870 ^ x163;
  assign n4872 = x752 ^ x703;
  assign n4873 = n4872 ^ x752;
  assign n4874 = x907 ^ x752;
  assign n4875 = n4874 ^ x752;
  assign n4876 = n4873 & n4875;
  assign n4877 = n4876 ^ x752;
  assign n4878 = ~x947 & ~n4877;
  assign n4879 = n4878 ^ x752;
  assign n4880 = n4879 ^ x164;
  assign n4881 = ~n4554 & n4880;
  assign n4882 = n4881 ^ x164;
  assign n4883 = x907 ^ x774;
  assign n4884 = n4883 ^ x774;
  assign n4885 = n4643 & n4884;
  assign n4886 = n4885 ^ x774;
  assign n4887 = ~x947 & ~n4886;
  assign n4888 = n4887 ^ x774;
  assign n4889 = ~n4710 & ~n4888;
  assign n4890 = ~x165 & n4554;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = x772 ^ x727;
  assign n4893 = n4892 ^ x772;
  assign n4894 = x907 ^ x772;
  assign n4895 = n4894 ^ x772;
  assign n4896 = n4893 & n4895;
  assign n4897 = n4896 ^ x772;
  assign n4898 = ~x947 & n4897;
  assign n4899 = n4898 ^ x772;
  assign n4900 = n4899 ^ x166;
  assign n4901 = ~n4554 & n4900;
  assign n4902 = n4901 ^ x166;
  assign n4903 = x768 ^ x705;
  assign n4904 = n4903 ^ x768;
  assign n4905 = x907 ^ x768;
  assign n4906 = n4905 ^ x768;
  assign n4907 = n4904 & n4906;
  assign n4908 = n4907 ^ x768;
  assign n4909 = ~x947 & ~n4908;
  assign n4910 = n4909 ^ x768;
  assign n4911 = n4910 ^ x167;
  assign n4912 = ~n4554 & n4911;
  assign n4913 = n4912 ^ x167;
  assign n4914 = x763 ^ x699;
  assign n4915 = n4914 ^ x763;
  assign n4916 = x907 ^ x763;
  assign n4917 = n4916 ^ x763;
  assign n4918 = n4915 & n4917;
  assign n4919 = n4918 ^ x763;
  assign n4920 = ~x947 & n4919;
  assign n4921 = n4920 ^ x763;
  assign n4922 = n4921 ^ x168;
  assign n4923 = ~n4554 & ~n4922;
  assign n4924 = n4923 ^ x168;
  assign n4925 = x746 ^ x729;
  assign n4926 = n4925 ^ x746;
  assign n4927 = x907 ^ x746;
  assign n4928 = n4927 ^ x746;
  assign n4929 = n4926 & n4928;
  assign n4930 = n4929 ^ x746;
  assign n4931 = ~x947 & n4930;
  assign n4932 = n4931 ^ x746;
  assign n4933 = n4932 ^ x169;
  assign n4934 = ~n4554 & ~n4933;
  assign n4935 = n4934 ^ x169;
  assign n4936 = x748 ^ x730;
  assign n4937 = n4936 ^ x748;
  assign n4938 = x907 ^ x748;
  assign n4939 = n4938 ^ x748;
  assign n4940 = n4937 & n4939;
  assign n4941 = n4940 ^ x748;
  assign n4942 = ~x947 & n4941;
  assign n4943 = n4942 ^ x748;
  assign n4944 = n4943 ^ x170;
  assign n4945 = ~n4554 & ~n4944;
  assign n4946 = n4945 ^ x170;
  assign n4947 = x764 ^ x691;
  assign n4948 = n4947 ^ x764;
  assign n4949 = x907 ^ x764;
  assign n4950 = n4949 ^ x764;
  assign n4951 = n4948 & n4950;
  assign n4952 = n4951 ^ x764;
  assign n4953 = ~x947 & n4952;
  assign n4954 = n4953 ^ x764;
  assign n4955 = n4954 ^ x171;
  assign n4956 = ~n4554 & ~n4955;
  assign n4957 = n4956 ^ x171;
  assign n4958 = x739 ^ x690;
  assign n4959 = n4958 ^ x739;
  assign n4960 = x907 ^ x739;
  assign n4961 = n4960 ^ x739;
  assign n4962 = n4959 & n4961;
  assign n4963 = n4962 ^ x739;
  assign n4964 = ~x947 & n4963;
  assign n4965 = n4964 ^ x739;
  assign n4966 = n4965 ^ x172;
  assign n4967 = ~n4554 & ~n4966;
  assign n4968 = n4967 ^ x172;
  assign n4969 = n4606 ^ x745;
  assign n4970 = n4969 ^ x745;
  assign n4971 = ~n4734 & n4970;
  assign n4972 = n4971 ^ x745;
  assign n4973 = ~n4580 & ~n4972;
  assign n4974 = n4973 ^ x745;
  assign n4975 = n4974 ^ x173;
  assign n4976 = ~n4554 & n4975;
  assign n4977 = n4976 ^ x173;
  assign n4978 = n4606 ^ x759;
  assign n4979 = n4978 ^ x759;
  assign n4980 = n4745 & n4979;
  assign n4981 = n4980 ^ x759;
  assign n4982 = ~n4580 & n4981;
  assign n4983 = n4982 ^ x759;
  assign n4984 = n4983 ^ x174;
  assign n4985 = ~n4554 & n4984;
  assign n4986 = n4985 ^ x174;
  assign n4987 = n4606 ^ x766;
  assign n4988 = n4987 ^ x766;
  assign n4989 = n4756 & n4988;
  assign n4990 = n4989 ^ x766;
  assign n4991 = ~n4580 & n4990;
  assign n4992 = n4991 ^ x766;
  assign n4993 = n4992 ^ x175;
  assign n4994 = ~n4554 & ~n4993;
  assign n4995 = n4994 ^ x175;
  assign n4996 = n4606 ^ x742;
  assign n4997 = n4996 ^ x742;
  assign n4998 = ~n4767 & n4997;
  assign n4999 = n4998 ^ x742;
  assign n5000 = ~n4580 & ~n4999;
  assign n5001 = n5000 ^ x742;
  assign n5002 = n5001 ^ x176;
  assign n5003 = ~n4554 & n5002;
  assign n5004 = n5003 ^ x176;
  assign n5005 = n4606 ^ x757;
  assign n5006 = n5005 ^ x757;
  assign n5007 = ~n4778 & n5006;
  assign n5008 = n5007 ^ x757;
  assign n5009 = ~n4580 & ~n5008;
  assign n5010 = n5009 ^ x757;
  assign n5011 = n5010 ^ x177;
  assign n5012 = ~n4554 & n5011;
  assign n5013 = n5012 ^ x177;
  assign n5014 = n4606 ^ x760;
  assign n5015 = n5014 ^ x760;
  assign n5016 = ~n4800 & n5015;
  assign n5017 = n5016 ^ x760;
  assign n5018 = ~n4580 & ~n5017;
  assign n5019 = n5018 ^ x760;
  assign n5020 = n5019 ^ x178;
  assign n5021 = ~n4554 & n5020;
  assign n5022 = n5021 ^ x178;
  assign n5023 = n4606 ^ x741;
  assign n5024 = n5023 ^ x741;
  assign n5025 = ~n4789 & n5024;
  assign n5026 = n5025 ^ x741;
  assign n5027 = ~n4580 & ~n5026;
  assign n5028 = n5027 ^ x741;
  assign n5029 = n5028 ^ x179;
  assign n5030 = ~n4554 & n5029;
  assign n5031 = n5030 ^ x179;
  assign n5032 = n4606 ^ x753;
  assign n5033 = n5032 ^ x753;
  assign n5034 = ~n4811 & n5033;
  assign n5035 = n5034 ^ x753;
  assign n5036 = ~n4580 & ~n5035;
  assign n5037 = n5036 ^ x753;
  assign n5038 = n5037 ^ x180;
  assign n5039 = ~n4554 & n5038;
  assign n5040 = n5039 ^ x180;
  assign n5041 = n4606 ^ x754;
  assign n5042 = n5041 ^ x754;
  assign n5043 = ~n4822 & n5042;
  assign n5044 = n5043 ^ x754;
  assign n5045 = ~n4580 & ~n5044;
  assign n5046 = n5045 ^ x754;
  assign n5047 = n5046 ^ x181;
  assign n5048 = ~n4554 & n5047;
  assign n5049 = n5048 ^ x181;
  assign n5050 = n4606 ^ x756;
  assign n5051 = n5050 ^ x756;
  assign n5052 = ~n4833 & n5051;
  assign n5053 = n5052 ^ x756;
  assign n5054 = ~n4580 & ~n5053;
  assign n5055 = n5054 ^ x756;
  assign n5056 = n5055 ^ x182;
  assign n5057 = ~n4554 & n5056;
  assign n5058 = n5057 ^ x182;
  assign n5059 = n4606 ^ x755;
  assign n5060 = n5059 ^ x755;
  assign n5061 = ~n4712 & n5060;
  assign n5062 = n5061 ^ x755;
  assign n5063 = ~n4580 & ~n5062;
  assign n5064 = n5063 ^ x755;
  assign n5065 = n5064 ^ x183;
  assign n5066 = ~n4554 & n5065;
  assign n5067 = n5066 ^ x183;
  assign n5068 = n4606 ^ x777;
  assign n5069 = n5068 ^ x777;
  assign n5070 = ~n4862 & n5069;
  assign n5071 = n5070 ^ x777;
  assign n5072 = ~n4580 & ~n5071;
  assign n5073 = n5072 ^ x777;
  assign n5074 = n5073 ^ x184;
  assign n5075 = ~n4554 & n5074;
  assign n5076 = n5075 ^ x184;
  assign n5077 = n4606 ^ x751;
  assign n5078 = n5077 ^ x751;
  assign n5079 = ~n4723 & n5078;
  assign n5080 = n5079 ^ x751;
  assign n5081 = ~n4580 & ~n5080;
  assign n5082 = n5081 ^ x751;
  assign n5083 = n5082 ^ x185;
  assign n5084 = ~n4554 & n5083;
  assign n5085 = n5084 ^ x185;
  assign n5086 = n4606 ^ x752;
  assign n5087 = n5086 ^ x752;
  assign n5088 = n4873 & n5087;
  assign n5089 = n5088 ^ x752;
  assign n5090 = ~n4580 & ~n5089;
  assign n5091 = n5090 ^ x752;
  assign n5092 = n5091 ^ x186;
  assign n5093 = ~n4554 & n5092;
  assign n5094 = n5093 ^ x186;
  assign n5095 = n4606 ^ x770;
  assign n5096 = n5095 ^ x770;
  assign n5097 = n4683 & n5096;
  assign n5098 = n5097 ^ x770;
  assign n5099 = ~n4580 & ~n5098;
  assign n5100 = n5099 ^ x770;
  assign n5101 = n5100 ^ x187;
  assign n5102 = ~n4554 & n5101;
  assign n5103 = n5102 ^ x187;
  assign n5104 = n4606 ^ x768;
  assign n5105 = n5104 ^ x768;
  assign n5106 = n4904 & n5105;
  assign n5107 = n5106 ^ x768;
  assign n5108 = ~n4580 & ~n5107;
  assign n5109 = n5108 ^ x768;
  assign n5110 = n5109 ^ x188;
  assign n5111 = ~n4554 & n5110;
  assign n5112 = n5111 ^ x188;
  assign n5113 = n4606 ^ x772;
  assign n5114 = n5113 ^ x772;
  assign n5115 = n4893 & n5114;
  assign n5116 = n5115 ^ x772;
  assign n5117 = ~n4580 & n5116;
  assign n5118 = n5117 ^ x772;
  assign n5119 = n5118 ^ x189;
  assign n5120 = ~n4554 & n5119;
  assign n5121 = n5120 ^ x189;
  assign n5122 = n4606 ^ x763;
  assign n5123 = n5122 ^ x763;
  assign n5124 = n4915 & n5123;
  assign n5125 = n5124 ^ x763;
  assign n5126 = ~n4580 & n5125;
  assign n5127 = n5126 ^ x763;
  assign n5128 = n5127 ^ x190;
  assign n5129 = ~n4554 & ~n5128;
  assign n5130 = n5129 ^ x190;
  assign n5131 = n4606 ^ x746;
  assign n5132 = n5131 ^ x746;
  assign n5133 = n4926 & n5132;
  assign n5134 = n5133 ^ x746;
  assign n5135 = ~n4580 & n5134;
  assign n5136 = n5135 ^ x746;
  assign n5137 = n5136 ^ x191;
  assign n5138 = ~n4554 & ~n5137;
  assign n5139 = n5138 ^ x191;
  assign n5140 = n4606 ^ x764;
  assign n5141 = n5140 ^ x764;
  assign n5142 = n4948 & n5141;
  assign n5143 = n5142 ^ x764;
  assign n5144 = ~n4580 & n5143;
  assign n5145 = n5144 ^ x764;
  assign n5146 = n5145 ^ x192;
  assign n5147 = ~n4554 & ~n5146;
  assign n5148 = n5147 ^ x192;
  assign n5149 = n4606 ^ x739;
  assign n5150 = n5149 ^ x739;
  assign n5151 = n4959 & n5150;
  assign n5152 = n5151 ^ x739;
  assign n5153 = ~n4580 & n5152;
  assign n5154 = n5153 ^ x739;
  assign n5155 = n5154 ^ x193;
  assign n5156 = ~n4554 & ~n5155;
  assign n5157 = n5156 ^ x193;
  assign n5158 = n4606 ^ x748;
  assign n5159 = n5158 ^ x748;
  assign n5160 = n4937 & n5159;
  assign n5161 = n5160 ^ x748;
  assign n5162 = ~n4580 & n5161;
  assign n5163 = n5162 ^ x748;
  assign n5164 = n5163 ^ x194;
  assign n5165 = ~n4554 & ~n5164;
  assign n5166 = n5165 ^ x194;
  assign n5167 = ~x299 & n4426;
  assign n5168 = n5167 ^ x171;
  assign n5169 = n2643 & n5168;
  assign n5170 = n5169 ^ n4513;
  assign n5171 = n5170 ^ n5169;
  assign n5172 = n2954 & n3980;
  assign n5173 = ~x196 & n5172;
  assign n5174 = x195 & ~n5173;
  assign n5175 = n5174 ^ n5169;
  assign n5176 = n5175 ^ n5169;
  assign n5177 = n5171 & n5176;
  assign n5178 = n5177 ^ n5169;
  assign n5179 = n3607 & ~n5178;
  assign n5180 = n5179 ^ n5169;
  assign n5181 = ~x299 & n4449;
  assign n5182 = n5181 ^ x170;
  assign n5183 = n2643 & n5182;
  assign n5184 = n5183 ^ n4513;
  assign n5185 = n5184 ^ n5183;
  assign n5187 = ~x195 & n5173;
  assign n5186 = n5172 ^ x196;
  assign n5188 = n5187 ^ n5186;
  assign n5189 = n5188 ^ n5183;
  assign n5190 = n5189 ^ n5183;
  assign n5191 = n5185 & n5190;
  assign n5192 = n5191 ^ n5183;
  assign n5193 = n3607 & ~n5192;
  assign n5194 = n5193 ^ n5183;
  assign n5195 = x907 ^ x767;
  assign n5196 = n5195 ^ x767;
  assign n5197 = ~n4665 & n5196;
  assign n5198 = n5197 ^ x767;
  assign n5199 = ~x947 & ~n5198;
  assign n5200 = n5199 ^ x767;
  assign n5201 = n5200 ^ x197;
  assign n5202 = ~n4554 & n5201;
  assign n5203 = n5202 ^ x197;
  assign n5204 = n4606 ^ x633;
  assign n5205 = n5204 ^ x633;
  assign n5206 = x634 ^ x633;
  assign n5207 = n5206 ^ x633;
  assign n5208 = n5205 & n5207;
  assign n5209 = n5208 ^ x633;
  assign n5210 = ~n4580 & n5209;
  assign n5211 = n5210 ^ x633;
  assign n5212 = n5211 ^ x198;
  assign n5213 = n4552 & n5212;
  assign n5214 = n5213 ^ x198;
  assign n5215 = n4606 ^ x617;
  assign n5216 = n5215 ^ x617;
  assign n5217 = x637 ^ x617;
  assign n5218 = n5217 ^ x617;
  assign n5219 = n5216 & n5218;
  assign n5220 = n5219 ^ x617;
  assign n5221 = ~n4580 & n5220;
  assign n5222 = n5221 ^ x617;
  assign n5223 = n5222 ^ x199;
  assign n5224 = n4552 & n5223;
  assign n5225 = n5224 ^ x199;
  assign n5226 = x643 ^ x606;
  assign n5227 = n5226 ^ x606;
  assign n5228 = n4606 ^ x606;
  assign n5229 = n5228 ^ x606;
  assign n5230 = n5227 & n5229;
  assign n5231 = n5230 ^ x606;
  assign n5232 = ~n4580 & n5231;
  assign n5233 = n5232 ^ x606;
  assign n5234 = n5233 ^ x200;
  assign n5235 = n4552 & n5234;
  assign n5236 = n5235 ^ x200;
  assign n5237 = ~n1241 & n3448;
  assign n5238 = ~x332 & ~n1601;
  assign n5239 = ~n5237 & n5238;
  assign n5241 = n1257 & ~n1729;
  assign n5242 = n5241 ^ x198;
  assign n5240 = ~x32 & x70;
  assign n5243 = n5242 ^ n5240;
  assign n5244 = n5240 ^ x96;
  assign n5245 = n5244 ^ x96;
  assign n5246 = ~x70 & n2921;
  assign n5247 = n5246 ^ x96;
  assign n5248 = ~n5245 & n5247;
  assign n5249 = n5248 ^ x96;
  assign n5250 = ~n5243 & ~n5249;
  assign n5251 = n5250 ^ n5242;
  assign n5252 = x233 & ~n5251;
  assign n5253 = x237 & n5252;
  assign n5254 = n5239 & ~n5253;
  assign n5255 = ~n2346 & n2349;
  assign n5256 = ~x587 & ~n5255;
  assign n5257 = n5256 ^ n2519;
  assign n5258 = n5256 ^ n2346;
  assign n5259 = n5256 ^ n1729;
  assign n5260 = ~n5256 & ~n5259;
  assign n5261 = n5260 ^ n5256;
  assign n5262 = n5258 & ~n5261;
  assign n5263 = n5262 ^ n5260;
  assign n5264 = n5263 ^ n5256;
  assign n5265 = n5264 ^ n1729;
  assign n5266 = ~n5257 & ~n5265;
  assign n5267 = n5266 ^ n2519;
  assign n5268 = ~x332 & ~n5267;
  assign n5269 = ~n5254 & ~n5268;
  assign n5270 = ~x201 & ~n5269;
  assign n5271 = x96 & n5242;
  assign n5272 = x237 & n5271;
  assign n5273 = x233 & n5267;
  assign n5274 = n5272 & n5273;
  assign n5275 = ~n5270 & ~n5274;
  assign n5276 = ~x233 & ~n5251;
  assign n5277 = x237 & n5276;
  assign n5278 = n5239 & ~n5277;
  assign n5279 = ~n5268 & ~n5278;
  assign n5280 = ~x202 & ~n5279;
  assign n5281 = ~x233 & n5267;
  assign n5282 = n5272 & n5281;
  assign n5283 = ~n5280 & ~n5282;
  assign n5284 = ~x237 & n5276;
  assign n5285 = n5239 & ~n5284;
  assign n5286 = ~n5268 & ~n5285;
  assign n5287 = ~x203 & ~n5286;
  assign n5288 = ~x237 & n5271;
  assign n5289 = n5281 & n5288;
  assign n5290 = ~n5287 & ~n5289;
  assign n5291 = n1729 ^ x907;
  assign n5292 = n5291 ^ x907;
  assign n5293 = x907 ^ x602;
  assign n5294 = n5292 & n5293;
  assign n5295 = n5294 ^ x907;
  assign n5296 = n5295 ^ n2352;
  assign n5297 = n2346 & n5296;
  assign n5298 = n5297 ^ n2352;
  assign n5299 = ~x332 & ~n5298;
  assign n5300 = ~n5254 & ~n5299;
  assign n5301 = ~x204 & ~n5300;
  assign n5302 = n5272 & n5298;
  assign n5303 = x233 & n5302;
  assign n5304 = ~n5301 & ~n5303;
  assign n5305 = ~n5278 & ~n5299;
  assign n5306 = ~x205 & ~n5305;
  assign n5307 = ~x233 & n5302;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = ~x237 & n5252;
  assign n5310 = n5239 & ~n5309;
  assign n5311 = ~n5299 & ~n5310;
  assign n5312 = ~x206 & ~n5311;
  assign n5313 = n5288 & n5298;
  assign n5314 = x233 & n5313;
  assign n5315 = ~n5312 & ~n5314;
  assign n5316 = n4606 ^ x623;
  assign n5317 = n5316 ^ x623;
  assign n5318 = x710 ^ x623;
  assign n5319 = n5318 ^ x623;
  assign n5320 = n5317 & n5319;
  assign n5321 = n5320 ^ x623;
  assign n5322 = ~n4580 & n5321;
  assign n5323 = n5322 ^ x623;
  assign n5324 = n5323 ^ x207;
  assign n5325 = n4552 & ~n5324;
  assign n5326 = n5325 ^ x207;
  assign n5327 = x638 ^ x607;
  assign n5328 = n5327 ^ x607;
  assign n5329 = n4606 ^ x607;
  assign n5330 = n5329 ^ x607;
  assign n5331 = n5328 & n5330;
  assign n5332 = n5331 ^ x607;
  assign n5333 = ~n4580 & n5332;
  assign n5334 = n5333 ^ x607;
  assign n5335 = n5334 ^ x208;
  assign n5336 = n4552 & ~n5335;
  assign n5337 = n5336 ^ x208;
  assign n5338 = x639 ^ x622;
  assign n5339 = n5338 ^ x622;
  assign n5340 = n4606 ^ x622;
  assign n5341 = n5340 ^ x622;
  assign n5342 = n5339 & n5341;
  assign n5343 = n5342 ^ x622;
  assign n5344 = ~n4580 & n5343;
  assign n5345 = n5344 ^ x622;
  assign n5346 = n5345 ^ x209;
  assign n5347 = n4552 & ~n5346;
  assign n5348 = n5347 ^ x209;
  assign n5349 = x907 ^ x633;
  assign n5350 = n5349 ^ x633;
  assign n5351 = n5207 & n5350;
  assign n5352 = n5351 ^ x633;
  assign n5353 = ~x947 & n5352;
  assign n5354 = n5353 ^ x633;
  assign n5355 = n5354 ^ x210;
  assign n5356 = n4552 & n5355;
  assign n5357 = n5356 ^ x210;
  assign n5358 = x907 ^ x606;
  assign n5359 = n5358 ^ x606;
  assign n5360 = n5227 & n5359;
  assign n5361 = n5360 ^ x606;
  assign n5362 = ~x947 & n5361;
  assign n5363 = n5362 ^ x606;
  assign n5364 = n5363 ^ x211;
  assign n5365 = n4552 & n5364;
  assign n5366 = n5365 ^ x211;
  assign n5367 = ~x212 & ~n4552;
  assign n5368 = x907 ^ x607;
  assign n5369 = n5368 ^ x607;
  assign n5370 = n5328 & n5369;
  assign n5371 = n5370 ^ x607;
  assign n5372 = ~x947 & n5371;
  assign n5373 = n5372 ^ x607;
  assign n5374 = n4709 & n5373;
  assign n5375 = ~n5367 & ~n5374;
  assign n5376 = ~x213 & ~n4552;
  assign n5377 = x907 ^ x622;
  assign n5378 = n5377 ^ x622;
  assign n5379 = n5339 & n5378;
  assign n5380 = n5379 ^ x622;
  assign n5381 = ~x947 & n5380;
  assign n5382 = n5381 ^ x622;
  assign n5383 = n4709 & n5382;
  assign n5384 = ~n5376 & ~n5383;
  assign n5385 = x907 ^ x623;
  assign n5386 = n5385 ^ x623;
  assign n5387 = n5319 & n5386;
  assign n5388 = n5387 ^ x623;
  assign n5389 = ~x947 & n5388;
  assign n5390 = n5389 ^ x623;
  assign n5391 = n5390 ^ x214;
  assign n5392 = n4552 & ~n5391;
  assign n5393 = n5392 ^ x214;
  assign n5394 = x681 ^ x642;
  assign n5395 = n5394 ^ x642;
  assign n5396 = x907 ^ x642;
  assign n5397 = n5396 ^ x642;
  assign n5398 = n5395 & n5397;
  assign n5399 = n5398 ^ x642;
  assign n5400 = ~x947 & n5399;
  assign n5401 = n5400 ^ x642;
  assign n5402 = n5401 ^ x215;
  assign n5403 = n4552 & n5402;
  assign n5404 = n5403 ^ x215;
  assign n5405 = x662 ^ x614;
  assign n5406 = n5405 ^ x614;
  assign n5407 = x907 ^ x614;
  assign n5408 = n5407 ^ x614;
  assign n5409 = n5406 & n5408;
  assign n5410 = n5409 ^ x614;
  assign n5411 = ~x947 & n5410;
  assign n5412 = n5411 ^ x614;
  assign n5413 = n5412 ^ x216;
  assign n5414 = n4552 & n5413;
  assign n5415 = n5414 ^ x216;
  assign n5416 = n4606 ^ x612;
  assign n5417 = n5416 ^ x612;
  assign n5418 = x695 ^ x612;
  assign n5419 = n5418 ^ x612;
  assign n5420 = n5417 & ~n5419;
  assign n5421 = n5420 ^ x612;
  assign n5422 = ~n4580 & n5421;
  assign n5423 = n5422 ^ x612;
  assign n5424 = n5423 ^ x217;
  assign n5425 = n4552 & ~n5424;
  assign n5426 = n5425 ^ x217;
  assign n5427 = ~n5285 & ~n5299;
  assign n5428 = ~x218 & ~n5427;
  assign n5429 = ~x233 & n5313;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431 = x219 & ~n4552;
  assign n5432 = x907 ^ x617;
  assign n5433 = n5432 ^ x617;
  assign n5434 = n5218 & n5433;
  assign n5435 = n5434 ^ x617;
  assign n5436 = ~x947 & n5435;
  assign n5437 = n5436 ^ x617;
  assign n5438 = n4709 & n5437;
  assign n5439 = ~n5431 & ~n5438;
  assign n5440 = ~n5268 & ~n5310;
  assign n5441 = ~x220 & ~n5440;
  assign n5442 = n5273 & n5288;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = x661 ^ x616;
  assign n5445 = n5444 ^ x616;
  assign n5446 = x907 ^ x616;
  assign n5447 = n5446 ^ x616;
  assign n5448 = n5445 & n5447;
  assign n5449 = n5448 ^ x616;
  assign n5450 = ~x947 & n5449;
  assign n5451 = n5450 ^ x616;
  assign n5452 = n5451 ^ x221;
  assign n5453 = n4552 & n5452;
  assign n5454 = n5453 ^ x221;
  assign n5455 = n4606 ^ x616;
  assign n5456 = n5455 ^ x616;
  assign n5457 = n5445 & n5456;
  assign n5458 = n5457 ^ x616;
  assign n5459 = ~n4580 & n5458;
  assign n5460 = n5459 ^ x616;
  assign n5461 = n5460 ^ x222;
  assign n5462 = n4552 & n5461;
  assign n5463 = n5462 ^ x222;
  assign n5464 = n4606 ^ x642;
  assign n5465 = n5464 ^ x642;
  assign n5466 = n5395 & n5465;
  assign n5467 = n5466 ^ x642;
  assign n5468 = ~n4580 & n5467;
  assign n5469 = n5468 ^ x642;
  assign n5470 = n5469 ^ x223;
  assign n5471 = n4552 & n5470;
  assign n5472 = n5471 ^ x223;
  assign n5473 = n4606 ^ x614;
  assign n5474 = n5473 ^ x614;
  assign n5475 = n5406 & n5474;
  assign n5476 = n5475 ^ x614;
  assign n5477 = ~n4580 & n5476;
  assign n5478 = n5477 ^ x614;
  assign n5479 = n5478 ^ x224;
  assign n5480 = n4552 & n5479;
  assign n5481 = n5480 ^ x224;
  assign n5482 = n1524 & n1572;
  assign n5483 = x70 & x332;
  assign n5484 = ~n1262 & ~n5483;
  assign n5485 = n1752 & ~n5484;
  assign n5486 = n1497 & n4044;
  assign n5487 = ~x55 & ~x137;
  assign n5488 = ~n5486 & n5487;
  assign n5489 = ~n1632 & ~n5488;
  assign n5490 = ~n5485 & ~n5489;
  assign n5491 = ~n5482 & n5490;
  assign n5492 = n1752 & n2311;
  assign n5493 = n1614 & ~n1619;
  assign n5494 = x479 & n3851;
  assign n5495 = n1631 & ~n5494;
  assign n5496 = ~n5493 & n5495;
  assign n5497 = ~n5492 & n5496;
  assign n5498 = n5497 ^ x231;
  assign n5499 = ~x228 & ~n5498;
  assign n5500 = n5499 ^ x231;
  assign n5501 = x1093 & n3259;
  assign n5502 = ~x58 & n1504;
  assign n5503 = n1308 & n5502;
  assign n5504 = ~x72 & ~n5503;
  assign n5505 = ~n3431 & n5504;
  assign n5506 = ~n5501 & n5505;
  assign n5507 = n1752 & ~n5506;
  assign n5508 = ~n3603 & ~n5507;
  assign n5509 = x36 & n1478;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = ~n1471 & ~n2319;
  assign n5512 = n1571 & n1658;
  assign n5513 = ~n5511 & n5512;
  assign n5514 = ~n1470 & n5513;
  assign n5515 = ~x228 & ~n5514;
  assign n5516 = ~x39 & ~n5515;
  assign n5517 = x1091 & n3843;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = ~x47 & ~n2320;
  assign n5520 = n1233 & n5519;
  assign n5521 = ~n2973 & n5520;
  assign n5522 = ~n4551 & ~n5521;
  assign n5523 = ~x64 & n2962;
  assign n5524 = x102 ^ x65;
  assign n5525 = n5523 & n5524;
  assign n5526 = n1398 & n5525;
  assign n5527 = ~n3218 & ~n5526;
  assign n5528 = ~n2414 & n5527;
  assign n5529 = ~n1632 & ~n3546;
  assign n5530 = ~n5528 & ~n5529;
  assign n5558 = ~x209 & n1729;
  assign n5533 = x208 ^ x207;
  assign n5559 = x199 & ~x200;
  assign n5560 = x1154 & n5559;
  assign n5561 = x1156 ^ x1155;
  assign n5562 = x1155 ^ x200;
  assign n5563 = n5562 ^ x1155;
  assign n5564 = n5561 & ~n5563;
  assign n5565 = n5564 ^ x1155;
  assign n5566 = ~x199 & n5565;
  assign n5567 = ~n5560 & ~n5566;
  assign n5568 = n5567 ^ x208;
  assign n5569 = n5568 ^ n5567;
  assign n5570 = x200 ^ x199;
  assign n5571 = n5561 & n5563;
  assign n5572 = n5571 ^ x1155;
  assign n5573 = n5572 ^ x200;
  assign n5574 = n5573 ^ n5572;
  assign n5575 = n5572 ^ x1157;
  assign n5576 = n5575 ^ n5572;
  assign n5577 = ~n5574 & n5576;
  assign n5578 = n5577 ^ n5572;
  assign n5579 = ~n5570 & n5578;
  assign n5580 = n5579 ^ n5572;
  assign n5581 = n5580 ^ n5567;
  assign n5582 = ~n5569 & ~n5581;
  assign n5583 = n5582 ^ n5567;
  assign n5584 = n5533 & ~n5583;
  assign n5585 = n5558 & ~n5584;
  assign n5586 = x1154 & n3481;
  assign n5587 = x1153 & n5559;
  assign n5588 = ~n5586 & ~n5587;
  assign n5589 = x1155 & n3378;
  assign n5590 = n5588 & ~n5589;
  assign n5591 = n3381 & ~n5590;
  assign n5592 = n5585 & ~n5591;
  assign n5593 = n5592 ^ x233;
  assign n5594 = n5593 ^ x233;
  assign n5531 = x1142 & ~n3378;
  assign n5532 = ~n3382 & n5531;
  assign n5534 = n5533 ^ x200;
  assign n5535 = n5534 ^ x1143;
  assign n5536 = n5535 ^ x1143;
  assign n5537 = n5536 ^ n5533;
  assign n5538 = n5537 ^ n5536;
  assign n5539 = x1144 & n5538;
  assign n5540 = n5539 ^ x1143;
  assign n5541 = x1143 ^ x208;
  assign n5542 = ~n5537 & ~n5541;
  assign n5543 = n5542 ^ n5536;
  assign n5544 = n5543 ^ n5537;
  assign n5545 = n5540 & n5544;
  assign n5546 = ~n5536 & n5545;
  assign n5547 = n5546 ^ n5539;
  assign n5548 = ~n5532 & ~n5547;
  assign n5549 = ~x207 & ~x208;
  assign n5550 = ~x200 & ~n5549;
  assign n5551 = x1142 & n5550;
  assign n5552 = x199 & ~n5551;
  assign n5553 = ~n5548 & ~n5552;
  assign n5554 = x209 & n1729;
  assign n5555 = ~n5553 & n5554;
  assign n5556 = n5555 ^ x233;
  assign n5557 = n5556 ^ x233;
  assign n5595 = n5594 ^ n5557;
  assign n5607 = x1154 ^ x214;
  assign n5608 = n5607 ^ x1154;
  assign n5609 = x1155 ^ x1154;
  assign n5610 = ~n5608 & n5609;
  assign n5611 = n5610 ^ x1154;
  assign n5596 = x1156 ^ x1154;
  assign n5597 = ~x219 & n5596;
  assign n5598 = n5597 ^ x1154;
  assign n5599 = n5598 ^ x214;
  assign n5600 = n5599 ^ n5598;
  assign n5601 = x1155 ^ x1153;
  assign n5602 = ~x219 & n5601;
  assign n5603 = n5602 ^ x1153;
  assign n5604 = n5603 ^ n5598;
  assign n5605 = n5600 & n5604;
  assign n5606 = n5605 ^ n5598;
  assign n5612 = n5611 ^ n5606;
  assign n5613 = n5612 ^ n5606;
  assign n5614 = n5606 ^ x219;
  assign n5615 = n5614 ^ n5606;
  assign n5616 = n5613 & ~n5615;
  assign n5617 = n5616 ^ n5606;
  assign n5618 = x211 & n5617;
  assign n5619 = n5618 ^ n5606;
  assign n5620 = x212 & n5619;
  assign n5621 = ~x213 & ~n1729;
  assign n5622 = ~x212 & x214;
  assign n5623 = ~x219 & x1156;
  assign n5624 = n5623 ^ x211;
  assign n5625 = n5624 ^ n5623;
  assign n5626 = x1157 ^ x1155;
  assign n5627 = ~x219 & n5626;
  assign n5628 = n5627 ^ x1155;
  assign n5629 = n5628 ^ n5623;
  assign n5630 = ~n5625 & n5629;
  assign n5631 = n5630 ^ n5623;
  assign n5632 = n5622 & n5631;
  assign n5633 = n5621 & ~n5632;
  assign n5634 = ~n5620 & n5633;
  assign n5635 = ~x212 & ~x214;
  assign n5636 = n3477 & ~n5635;
  assign n5637 = x1143 & n5636;
  assign n5638 = n3384 & n3478;
  assign n5639 = n3475 & ~n5635;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = x1142 & ~n5640;
  assign n5642 = x214 ^ x212;
  assign n5643 = n3404 & n5642;
  assign n5644 = x1144 & n5643;
  assign n5645 = ~n5641 & ~n5644;
  assign n5646 = ~n5637 & n5645;
  assign n5647 = x213 & ~n1729;
  assign n5648 = n5646 & n5647;
  assign n5649 = ~n5634 & ~n5648;
  assign n5650 = n5649 ^ x233;
  assign n5651 = n5650 ^ x233;
  assign n5652 = n5651 ^ n5557;
  assign n5653 = ~n5557 & ~n5652;
  assign n5654 = n5653 ^ n5557;
  assign n5655 = n5595 & ~n5654;
  assign n5656 = n5655 ^ n5653;
  assign n5657 = n5656 ^ x233;
  assign n5658 = n5657 ^ n5557;
  assign n5659 = x230 & n5658;
  assign n5660 = n5659 ^ x233;
  assign n5661 = n5635 ^ n5549;
  assign n5662 = ~n1729 & n5661;
  assign n5663 = n5662 ^ n5549;
  assign n5664 = n3486 & ~n5663;
  assign n5665 = n3395 & n5664;
  assign n5666 = x1154 & n5665;
  assign n5667 = x1155 & n5636;
  assign n5668 = x1156 & n5643;
  assign n5669 = n5647 & ~n5668;
  assign n5670 = ~n5667 & n5669;
  assign n5671 = n5589 ^ n5566;
  assign n5672 = n5671 ^ n5566;
  assign n5673 = n5566 ^ x208;
  assign n5674 = n5673 ^ n5566;
  assign n5675 = n5672 & n5674;
  assign n5676 = n5675 ^ n5566;
  assign n5677 = ~n5533 & n5676;
  assign n5678 = n5677 ^ n5566;
  assign n5679 = n5554 & ~n5678;
  assign n5680 = ~n5670 & ~n5679;
  assign n5681 = ~n5666 & ~n5680;
  assign n5682 = n5681 ^ x234;
  assign n5683 = n5682 ^ x234;
  assign n5684 = x1152 & n5665;
  assign n5685 = ~n3395 & ~n5663;
  assign n5686 = x1154 ^ x1153;
  assign n5687 = n3486 ^ x1154;
  assign n5688 = n5687 ^ x1154;
  assign n5689 = n5686 & n5688;
  assign n5690 = n5689 ^ x1154;
  assign n5691 = n5685 & n5690;
  assign n5692 = ~n5684 & ~n5691;
  assign n5693 = ~n5554 & ~n5647;
  assign n5694 = n5692 & n5693;
  assign n5695 = n5694 ^ x234;
  assign n5696 = n5695 ^ x234;
  assign n5697 = ~n5683 & ~n5696;
  assign n5698 = n5697 ^ x234;
  assign n5699 = x230 & n5698;
  assign n5700 = n5699 ^ x234;
  assign n5701 = x213 & n5596;
  assign n5702 = n5701 ^ x1154;
  assign n5703 = n5636 & n5702;
  assign n5704 = x213 & n5601;
  assign n5705 = n5704 ^ x1153;
  assign n5706 = n5638 & n5705;
  assign n5707 = ~n1729 & ~n5706;
  assign n5708 = ~x211 & n5642;
  assign n5709 = n5603 ^ x213;
  assign n5710 = n5709 ^ n5603;
  assign n5711 = n5628 ^ n5603;
  assign n5712 = n5710 & n5711;
  assign n5713 = n5712 ^ n5603;
  assign n5714 = n5708 & n5713;
  assign n5715 = n5707 & ~n5714;
  assign n5716 = ~n5703 & n5715;
  assign n5717 = n5716 ^ x235;
  assign n5718 = n5717 ^ x235;
  assign n5719 = n5590 ^ n5580;
  assign n5720 = ~x209 & ~n5719;
  assign n5721 = n5720 ^ n5580;
  assign n5722 = n5533 & n5721;
  assign n5723 = x1153 ^ x200;
  assign n5724 = n5723 ^ x1153;
  assign n5725 = n5686 & ~n5724;
  assign n5726 = n5725 ^ x1153;
  assign n5727 = ~x199 & n5726;
  assign n5728 = n5558 & ~n5727;
  assign n5729 = x209 & ~n5566;
  assign n5730 = n3381 & ~n5729;
  assign n5731 = n1729 & ~n5730;
  assign n5732 = ~n5728 & ~n5731;
  assign n5733 = ~n5722 & ~n5732;
  assign n5734 = n5733 ^ x235;
  assign n5735 = n5734 ^ x235;
  assign n5736 = ~n5718 & ~n5735;
  assign n5737 = n5736 ^ x235;
  assign n5738 = x230 & n5737;
  assign n5739 = n5738 ^ x235;
  assign n5755 = x219 ^ x211;
  assign n5756 = x1156 ^ x219;
  assign n5757 = n5756 ^ x1156;
  assign n5758 = x1157 ^ x1156;
  assign n5759 = ~n5757 & n5758;
  assign n5760 = n5759 ^ x1156;
  assign n5761 = n5760 ^ x219;
  assign n5762 = n5761 ^ n5760;
  assign n5763 = n5760 ^ x1158;
  assign n5764 = n5763 ^ n5760;
  assign n5765 = ~n5762 & n5764;
  assign n5766 = n5765 ^ n5760;
  assign n5767 = ~n5755 & n5766;
  assign n5768 = n5767 ^ n5760;
  assign n5744 = n5628 ^ n5598;
  assign n5745 = ~x214 & n5744;
  assign n5746 = n5745 ^ n5598;
  assign n5740 = x1155 ^ x214;
  assign n5741 = n5740 ^ x1155;
  assign n5742 = n5561 & ~n5741;
  assign n5743 = n5742 ^ x1155;
  assign n5747 = n5746 ^ n5743;
  assign n5748 = n5747 ^ n5746;
  assign n5749 = n5746 ^ x219;
  assign n5750 = n5749 ^ n5746;
  assign n5751 = n5748 & ~n5750;
  assign n5752 = n5751 ^ n5746;
  assign n5753 = x211 & n5752;
  assign n5754 = n5753 ^ n5746;
  assign n5769 = n5768 ^ n5754;
  assign n5770 = n5769 ^ n5754;
  assign n5771 = n5754 ^ x214;
  assign n5772 = n5771 ^ n5754;
  assign n5773 = n5770 & n5772;
  assign n5774 = n5773 ^ n5754;
  assign n5775 = ~x212 & n5774;
  assign n5776 = n5775 ^ n5754;
  assign n5777 = n5621 & n5776;
  assign n5778 = n5580 ^ x208;
  assign n5779 = n5778 ^ n5580;
  assign n5780 = x1156 ^ x200;
  assign n5781 = n5780 ^ x1156;
  assign n5782 = n5758 & n5781;
  assign n5783 = n5782 ^ x1156;
  assign n5784 = n5783 ^ x200;
  assign n5785 = n5784 ^ n5783;
  assign n5786 = n5783 ^ x1158;
  assign n5787 = n5786 ^ n5783;
  assign n5788 = ~n5785 & n5787;
  assign n5789 = n5788 ^ n5783;
  assign n5790 = ~n5570 & n5789;
  assign n5791 = n5790 ^ n5783;
  assign n5792 = n5791 ^ n5580;
  assign n5793 = ~n5779 & n5792;
  assign n5794 = n5793 ^ n5580;
  assign n5795 = n5794 ^ x208;
  assign n5796 = n5795 ^ n5794;
  assign n5797 = n5794 ^ n5567;
  assign n5798 = n5797 ^ n5794;
  assign n5799 = n5796 & ~n5798;
  assign n5800 = n5799 ^ n5794;
  assign n5801 = ~n5533 & n5800;
  assign n5802 = n5801 ^ n5794;
  assign n5803 = n5558 & n5802;
  assign n5804 = x1143 & ~n5640;
  assign n5805 = ~x219 & n5642;
  assign n5806 = x1145 ^ x1144;
  assign n5807 = ~x211 & n5806;
  assign n5808 = n5807 ^ x1144;
  assign n5809 = n5805 & n5808;
  assign n5810 = n3384 & n3404;
  assign n5811 = x1144 & n5810;
  assign n5812 = ~n5809 & ~n5811;
  assign n5813 = ~n5804 & n5812;
  assign n5814 = n5647 & ~n5813;
  assign n5815 = x230 & ~n5814;
  assign n5816 = ~n5803 & n5815;
  assign n5817 = ~n5777 & n5816;
  assign n5818 = n5533 ^ n3381;
  assign n5819 = x200 & n5818;
  assign n5820 = n5819 ^ n3381;
  assign n5821 = x1144 & n5820;
  assign n5822 = x200 & x1143;
  assign n5823 = n3381 & n5822;
  assign n5824 = ~n5821 & ~n5823;
  assign n5825 = ~x199 & ~n5824;
  assign n5826 = n3381 ^ x1143;
  assign n5827 = n5826 ^ x1143;
  assign n5828 = x1145 ^ x1143;
  assign n5829 = n5828 ^ x1143;
  assign n5830 = ~n5827 & n5829;
  assign n5831 = n5830 ^ x1143;
  assign n5832 = ~x199 & n5831;
  assign n5833 = n5832 ^ x1143;
  assign n5834 = n5550 & n5833;
  assign n5835 = ~n5825 & ~n5834;
  assign n5836 = n5554 & ~n5835;
  assign n5837 = n5817 & ~n5836;
  assign n5838 = ~x230 & x237;
  assign n5839 = ~n5837 & ~n5838;
  assign n5848 = x1151 & n5665;
  assign n5849 = n3486 ^ x1153;
  assign n5850 = n5849 ^ x1153;
  assign n5851 = x1153 ^ x1152;
  assign n5852 = n5850 & n5851;
  assign n5853 = n5852 ^ x1153;
  assign n5854 = n5685 & n5853;
  assign n5855 = ~n5848 & ~n5854;
  assign n5856 = n5693 & n5855;
  assign n5857 = n5856 ^ x238;
  assign n5858 = n5857 ^ x238;
  assign n5840 = n3381 & ~n5587;
  assign n5841 = ~n5549 & ~n5840;
  assign n5842 = ~n5590 & n5841;
  assign n5843 = n5554 & ~n5842;
  assign n5844 = n3381 & n5727;
  assign n5845 = n5843 & ~n5844;
  assign n5846 = n5845 ^ x238;
  assign n5847 = n5846 ^ x238;
  assign n5859 = n5858 ^ n5847;
  assign n5860 = x1153 & ~n5640;
  assign n5861 = x1154 & n5810;
  assign n5862 = ~x211 & n5609;
  assign n5863 = n5862 ^ x1154;
  assign n5864 = n5805 & n5863;
  assign n5865 = ~n5861 & ~n5864;
  assign n5866 = ~n5860 & n5865;
  assign n5867 = n5647 & n5866;
  assign n5868 = n5867 ^ x238;
  assign n5869 = n5868 ^ x238;
  assign n5870 = n5869 ^ n5847;
  assign n5871 = ~n5847 & n5870;
  assign n5872 = n5871 ^ n5847;
  assign n5873 = n5859 & ~n5872;
  assign n5874 = n5873 ^ n5871;
  assign n5875 = n5874 ^ x238;
  assign n5876 = n5875 ^ n5847;
  assign n5877 = x230 & ~n5876;
  assign n5878 = n5877 ^ x238;
  assign n5879 = x207 & ~x208;
  assign n5880 = n1729 & n5879;
  assign n5881 = n5791 ^ n5567;
  assign n5882 = x209 & ~n5881;
  assign n5883 = n5882 ^ n5567;
  assign n5884 = n5880 & ~n5883;
  assign n5885 = n5884 ^ x239;
  assign n5886 = n5885 ^ x239;
  assign n5887 = ~n1729 & n5622;
  assign n5888 = n5754 ^ x213;
  assign n5889 = n5888 ^ n5754;
  assign n5890 = n5769 & n5889;
  assign n5891 = n5890 ^ n5754;
  assign n5892 = n5887 & n5891;
  assign n5893 = n5892 ^ x239;
  assign n5894 = n5893 ^ x239;
  assign n5895 = ~n5886 & ~n5894;
  assign n5896 = n5895 ^ x239;
  assign n5897 = x230 & ~n5896;
  assign n5898 = n5897 ^ x239;
  assign n5907 = x1147 & n5665;
  assign n5908 = n3486 ^ x1149;
  assign n5909 = n5908 ^ x1149;
  assign n5910 = x1149 ^ x1148;
  assign n5911 = n5909 & n5910;
  assign n5912 = n5911 ^ x1149;
  assign n5913 = n5685 & n5912;
  assign n5914 = ~n5907 & ~n5913;
  assign n5899 = x1145 & n5665;
  assign n5900 = n3486 ^ x1147;
  assign n5901 = n5900 ^ x1147;
  assign n5902 = x1147 ^ x1146;
  assign n5903 = n5901 & n5902;
  assign n5904 = n5903 ^ x1147;
  assign n5905 = n5685 & n5904;
  assign n5906 = ~n5899 & ~n5905;
  assign n5915 = n5914 ^ n5906;
  assign n5916 = ~n5693 & n5915;
  assign n5917 = n5916 ^ n5906;
  assign n5918 = n5917 ^ x240;
  assign n5919 = x230 & ~n5918;
  assign n5920 = n5919 ^ x240;
  assign n5921 = x1149 & n5665;
  assign n5922 = n3486 ^ x1151;
  assign n5923 = n5922 ^ x1151;
  assign n5924 = x1151 ^ x1150;
  assign n5925 = n5923 & n5924;
  assign n5926 = n5925 ^ x1151;
  assign n5927 = n5685 & n5926;
  assign n5928 = ~n5921 & ~n5927;
  assign n5929 = n5928 ^ n5855;
  assign n5930 = n5693 & n5929;
  assign n5931 = n5930 ^ n5855;
  assign n5932 = n5931 ^ x241;
  assign n5933 = x230 & ~n5932;
  assign n5934 = n5933 ^ x241;
  assign n5938 = x1144 & n5665;
  assign n5939 = n3486 ^ x1146;
  assign n5940 = n5939 ^ x1146;
  assign n5941 = x1146 ^ x1145;
  assign n5942 = n5940 & n5941;
  assign n5943 = n5942 ^ x1146;
  assign n5944 = n5685 & n5943;
  assign n5945 = ~n5938 & ~n5944;
  assign n5946 = ~n5693 & n5945;
  assign n5947 = n5946 ^ x242;
  assign n5948 = n5947 ^ x242;
  assign n5935 = n5621 & n5646;
  assign n5936 = n5935 ^ x242;
  assign n5937 = n5936 ^ x242;
  assign n5949 = n5948 ^ n5937;
  assign n5950 = ~n5553 & n5558;
  assign n5951 = n5950 ^ x242;
  assign n5952 = n5951 ^ x242;
  assign n5953 = n5952 ^ n5937;
  assign n5954 = ~n5937 & n5953;
  assign n5955 = n5954 ^ n5937;
  assign n5956 = n5949 & ~n5955;
  assign n5957 = n5956 ^ n5954;
  assign n5958 = n5957 ^ x242;
  assign n5959 = n5958 ^ n5937;
  assign n5960 = x230 & ~n5959;
  assign n5961 = n5960 ^ x242;
  assign n5962 = ~x230 & ~x1091;
  assign n5984 = n5559 ^ n3475;
  assign n5985 = n1729 & n5984;
  assign n5986 = n5985 ^ n3475;
  assign n5987 = x1157 & n5986;
  assign n5988 = ~n1729 & ~n3404;
  assign n5989 = ~n3380 & ~n5988;
  assign n5990 = x1155 & n5989;
  assign n5991 = ~n5987 & ~n5990;
  assign n5992 = ~n1729 & ~n3478;
  assign n5993 = ~n3483 & ~n5992;
  assign n5994 = x1156 & n5993;
  assign n5995 = n5991 & ~n5994;
  assign n5963 = ~x83 & ~x85;
  assign n5964 = n1729 ^ x199;
  assign n5965 = n5964 ^ x199;
  assign n5966 = n3552 & ~n5965;
  assign n5967 = n5966 ^ x199;
  assign n5968 = x81 & ~n5967;
  assign n5969 = n5963 & ~n5968;
  assign n5970 = x314 & ~n5969;
  assign n5971 = x802 & n5970;
  assign n5972 = x276 & n5971;
  assign n5973 = x271 & n5972;
  assign n5974 = x273 & n5973;
  assign n5975 = x283 & n5974;
  assign n5976 = x272 & n5975;
  assign n5977 = x275 & n5976;
  assign n5978 = x268 & n5977;
  assign n5979 = x253 & n5978;
  assign n5980 = x254 & n5979;
  assign n5981 = x267 & n5980;
  assign n5982 = ~x263 & n5981;
  assign n5983 = n5982 ^ x243;
  assign n5996 = n5995 ^ n5983;
  assign n5997 = ~n5962 & n5996;
  assign n5998 = n5997 ^ n5983;
  assign n6002 = ~n5693 & n5906;
  assign n6003 = n6002 ^ x244;
  assign n6004 = n6003 ^ x244;
  assign n5999 = n5558 & n5835;
  assign n6000 = n5999 ^ x244;
  assign n6001 = n6000 ^ x244;
  assign n6005 = n6004 ^ n6001;
  assign n6006 = n5621 & n5813;
  assign n6007 = n6006 ^ x244;
  assign n6008 = n6007 ^ x244;
  assign n6009 = n6008 ^ n6001;
  assign n6010 = ~n6001 & n6009;
  assign n6011 = n6010 ^ n6001;
  assign n6012 = n6005 & ~n6011;
  assign n6013 = n6012 ^ n6010;
  assign n6014 = n6013 ^ x244;
  assign n6015 = n6014 ^ n6001;
  assign n6016 = x230 & ~n6015;
  assign n6017 = n6016 ^ x244;
  assign n6018 = x1146 & n5665;
  assign n6019 = n3486 ^ x1148;
  assign n6020 = n6019 ^ x1148;
  assign n6021 = x1148 ^ x1147;
  assign n6022 = n6020 & n6021;
  assign n6023 = n6022 ^ x1148;
  assign n6024 = n5685 & n6023;
  assign n6025 = ~n6018 & ~n6024;
  assign n6026 = n6025 ^ n5945;
  assign n6027 = ~n5693 & n6026;
  assign n6028 = n6027 ^ n5945;
  assign n6029 = n6028 ^ x245;
  assign n6030 = x230 & ~n6029;
  assign n6031 = n6030 ^ x245;
  assign n6032 = x1148 & n5665;
  assign n6033 = n3486 ^ x1150;
  assign n6034 = n6033 ^ x1150;
  assign n6035 = x1150 ^ x1149;
  assign n6036 = n6034 & n6035;
  assign n6037 = n6036 ^ x1150;
  assign n6038 = n5685 & n6037;
  assign n6039 = ~n6032 & ~n6038;
  assign n6040 = n6039 ^ n6025;
  assign n6041 = ~n5693 & n6040;
  assign n6042 = n6041 ^ n6025;
  assign n6043 = n6042 ^ x246;
  assign n6044 = x230 & ~n6043;
  assign n6045 = n6044 ^ x246;
  assign n6046 = n5928 ^ n5914;
  assign n6047 = ~n5693 & n6046;
  assign n6048 = n6047 ^ n5914;
  assign n6049 = n6048 ^ x247;
  assign n6050 = x230 & ~n6049;
  assign n6051 = n6050 ^ x247;
  assign n6052 = x1150 & n5665;
  assign n6053 = n3486 ^ x1152;
  assign n6054 = n6053 ^ x1152;
  assign n6055 = x1152 ^ x1151;
  assign n6056 = n6054 & n6055;
  assign n6057 = n6056 ^ x1152;
  assign n6058 = n5685 & n6057;
  assign n6059 = ~n6052 & ~n6058;
  assign n6060 = n6059 ^ n6039;
  assign n6061 = ~n5693 & n6060;
  assign n6062 = n6061 ^ n6039;
  assign n6063 = n6062 ^ x248;
  assign n6064 = x230 & ~n6063;
  assign n6065 = n6064 ^ x248;
  assign n6066 = n6059 ^ n5692;
  assign n6067 = n5693 & n6066;
  assign n6068 = n6067 ^ n5692;
  assign n6069 = n6068 ^ x249;
  assign n6070 = x230 & ~n6069;
  assign n6071 = n6070 ^ x249;
  assign n6072 = ~n3460 & ~n4044;
  assign n6073 = ~x250 & ~n6072;
  assign n6074 = x1053 ^ x1039;
  assign n6075 = ~x200 & n6074;
  assign n6076 = n6075 ^ x1039;
  assign n6077 = n6076 ^ x251;
  assign n6078 = x476 ^ x200;
  assign n6079 = n6078 ^ x476;
  assign n6080 = x897 ^ x476;
  assign n6081 = ~n6079 & ~n6080;
  assign n6082 = n6081 ^ x476;
  assign n6083 = ~x199 & ~n6082;
  assign n6084 = n6077 & n6083;
  assign n6085 = n6084 ^ x251;
  assign n6086 = n2392 & ~n2396;
  assign n6087 = n2567 & n6086;
  assign n6088 = x1093 & ~n2872;
  assign n6089 = x252 & x1092;
  assign n6090 = ~n6088 & n6089;
  assign n6091 = ~n6087 & ~n6090;
  assign n6093 = x1153 & n5986;
  assign n6094 = x1151 & n5989;
  assign n6095 = ~n6093 & ~n6094;
  assign n6096 = x1152 & n5993;
  assign n6097 = n6095 & ~n6096;
  assign n6092 = n5978 ^ x253;
  assign n6098 = n6097 ^ n6092;
  assign n6099 = ~n5962 & ~n6098;
  assign n6100 = n6099 ^ n6092;
  assign n6102 = x1153 & n5993;
  assign n6103 = x1152 & n5989;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = x1154 & n5986;
  assign n6106 = n6104 & ~n6105;
  assign n6101 = n5979 ^ x254;
  assign n6107 = n6106 ^ n6101;
  assign n6108 = ~n5962 & ~n6107;
  assign n6109 = n6108 ^ n6101;
  assign n6110 = x1049 ^ x1036;
  assign n6111 = ~x200 & n6110;
  assign n6112 = n6111 ^ x1036;
  assign n6113 = n6112 ^ x255;
  assign n6114 = n6083 & n6113;
  assign n6115 = n6114 ^ x255;
  assign n6116 = x1070 ^ x1048;
  assign n6117 = x200 & n6116;
  assign n6118 = n6117 ^ x1048;
  assign n6119 = n6118 ^ x256;
  assign n6120 = n6083 & n6119;
  assign n6121 = n6120 ^ x256;
  assign n6122 = x1084 ^ x1065;
  assign n6123 = ~x200 & n6122;
  assign n6124 = n6123 ^ x1065;
  assign n6125 = n6124 ^ x257;
  assign n6126 = n6083 & n6125;
  assign n6127 = n6126 ^ x257;
  assign n6128 = x1072 ^ x1062;
  assign n6129 = ~x200 & n6128;
  assign n6130 = n6129 ^ x1062;
  assign n6131 = n6130 ^ x258;
  assign n6132 = n6083 & n6131;
  assign n6133 = n6132 ^ x258;
  assign n6134 = x1069 ^ x1059;
  assign n6135 = x200 & n6134;
  assign n6136 = n6135 ^ x1059;
  assign n6137 = n6136 ^ x259;
  assign n6138 = n6083 & n6137;
  assign n6139 = n6138 ^ x259;
  assign n6140 = x1067 ^ x1044;
  assign n6141 = x200 & n6140;
  assign n6142 = n6141 ^ x1044;
  assign n6143 = n6142 ^ x260;
  assign n6144 = n6083 & n6143;
  assign n6145 = n6144 ^ x260;
  assign n6146 = x1040 ^ x1037;
  assign n6147 = x200 & n6146;
  assign n6148 = n6147 ^ x1037;
  assign n6149 = n6148 ^ x261;
  assign n6150 = n6083 & n6149;
  assign n6151 = n6150 ^ x261;
  assign n6152 = x1093 ^ x123;
  assign n6153 = ~x228 & ~n6152;
  assign n6154 = n6153 ^ x123;
  assign n6155 = x1142 ^ x262;
  assign n6156 = n6155 ^ x262;
  assign n6157 = n5685 ^ x262;
  assign n6158 = n6157 ^ x262;
  assign n6159 = n6156 & n6158;
  assign n6160 = n6159 ^ x262;
  assign n6161 = ~n6154 & ~n6160;
  assign n6162 = n6161 ^ x262;
  assign n6164 = x1156 & n5986;
  assign n6165 = x1154 & n5989;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = x1155 & n5993;
  assign n6168 = n6166 & ~n6167;
  assign n6163 = n5981 ^ x263;
  assign n6169 = n6168 ^ n6163;
  assign n6170 = ~n5962 & n6169;
  assign n6171 = n6170 ^ n6163;
  assign n6177 = x796 ^ x264;
  assign n6178 = n5970 & ~n6177;
  assign n6179 = n6178 ^ x264;
  assign n6172 = x1141 & n5989;
  assign n6173 = x1143 & n5986;
  assign n6174 = ~n6172 & ~n6173;
  assign n6175 = x1142 & n5993;
  assign n6176 = n6174 & ~n6175;
  assign n6180 = n6179 ^ n6176;
  assign n6181 = ~n5962 & n6180;
  assign n6182 = n6181 ^ n6179;
  assign n6188 = x819 ^ x265;
  assign n6189 = n5970 & ~n6188;
  assign n6190 = n6189 ^ x265;
  assign n6183 = x1142 & n5989;
  assign n6184 = x1144 & n5986;
  assign n6185 = ~n6183 & ~n6184;
  assign n6186 = x1143 & n5993;
  assign n6187 = n6185 & ~n6186;
  assign n6191 = n6190 ^ n6187;
  assign n6192 = ~n5962 & n6191;
  assign n6193 = n6192 ^ n6190;
  assign n6199 = x948 ^ x266;
  assign n6200 = n5970 & n6199;
  assign n6201 = n6200 ^ x266;
  assign n6194 = x1134 & n5989;
  assign n6195 = x1136 & n5986;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = x1135 & n5993;
  assign n6198 = n6196 & ~n6197;
  assign n6202 = n6201 ^ n6198;
  assign n6203 = ~n5962 & ~n6202;
  assign n6204 = n6203 ^ n6201;
  assign n6206 = x1154 & n5993;
  assign n6207 = x1153 & n5989;
  assign n6208 = ~n6206 & ~n6207;
  assign n6209 = x1155 & n5986;
  assign n6210 = n6208 & ~n6209;
  assign n6205 = n5980 ^ x267;
  assign n6211 = n6210 ^ n6205;
  assign n6212 = ~n5962 & ~n6211;
  assign n6213 = n6212 ^ n6205;
  assign n6215 = x1152 & n5986;
  assign n6216 = x1150 & n5989;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = x1151 & n5993;
  assign n6219 = n6217 & ~n6218;
  assign n6214 = n5977 ^ x268;
  assign n6220 = n6219 ^ n6214;
  assign n6221 = ~n5962 & ~n6220;
  assign n6222 = n6221 ^ n6214;
  assign n6228 = x817 ^ x269;
  assign n6229 = n5970 & ~n6228;
  assign n6230 = n6229 ^ x269;
  assign n6223 = x1136 & n5989;
  assign n6224 = x1138 & n5986;
  assign n6225 = ~n6223 & ~n6224;
  assign n6226 = x1137 & n5993;
  assign n6227 = n6225 & ~n6226;
  assign n6231 = n6230 ^ n6227;
  assign n6232 = ~n5962 & n6231;
  assign n6233 = n6232 ^ n6230;
  assign n6239 = x805 ^ x270;
  assign n6240 = n5970 & ~n6239;
  assign n6241 = n6240 ^ x270;
  assign n6234 = x1139 & n5989;
  assign n6235 = x1141 & n5986;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = x1140 & n5993;
  assign n6238 = n6236 & ~n6237;
  assign n6242 = n6241 ^ n6238;
  assign n6243 = ~n5962 & n6242;
  assign n6244 = n6243 ^ n6241;
  assign n6246 = x1146 & n5993;
  assign n6247 = x1145 & n5989;
  assign n6248 = ~n6246 & ~n6247;
  assign n6249 = x1147 & n5986;
  assign n6250 = n6248 & ~n6249;
  assign n6245 = n5972 ^ x271;
  assign n6251 = n6250 ^ n6245;
  assign n6252 = ~n5962 & ~n6251;
  assign n6253 = n6252 ^ n6245;
  assign n6255 = x1150 & n5986;
  assign n6256 = x1148 & n5989;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = x1149 & n5993;
  assign n6259 = n6257 & ~n6258;
  assign n6254 = n5975 ^ x272;
  assign n6260 = n6259 ^ n6254;
  assign n6261 = ~n5962 & ~n6260;
  assign n6262 = n6261 ^ n6254;
  assign n6264 = x1146 & n5989;
  assign n6265 = x1148 & n5986;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = x1147 & n5993;
  assign n6268 = n6266 & ~n6267;
  assign n6263 = n5973 ^ x273;
  assign n6269 = n6268 ^ n6263;
  assign n6270 = ~n5962 & ~n6269;
  assign n6271 = n6270 ^ n6263;
  assign n6277 = x659 ^ x274;
  assign n6278 = n5970 & ~n6277;
  assign n6279 = n6278 ^ x274;
  assign n6272 = x1145 & n5986;
  assign n6273 = x1143 & n5989;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = x1144 & n5993;
  assign n6276 = n6274 & ~n6275;
  assign n6280 = n6279 ^ n6276;
  assign n6281 = ~n5962 & n6280;
  assign n6282 = n6281 ^ n6279;
  assign n6284 = x1151 & n5986;
  assign n6285 = x1149 & n5989;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = x1150 & n5993;
  assign n6288 = n6286 & ~n6287;
  assign n6283 = n5976 ^ x275;
  assign n6289 = n6288 ^ n6283;
  assign n6290 = ~n5962 & ~n6289;
  assign n6291 = n6290 ^ n6283;
  assign n6293 = x1146 & n5986;
  assign n6294 = x1144 & n5989;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = x1145 & n5993;
  assign n6297 = n6295 & ~n6296;
  assign n6292 = n5971 ^ x276;
  assign n6298 = n6297 ^ n6292;
  assign n6299 = ~n5962 & ~n6298;
  assign n6300 = n6299 ^ n6292;
  assign n6306 = x820 ^ x277;
  assign n6307 = n5970 & ~n6306;
  assign n6308 = n6307 ^ x277;
  assign n6301 = x1140 & n5989;
  assign n6302 = x1142 & n5986;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = x1141 & n5993;
  assign n6305 = n6303 & ~n6304;
  assign n6309 = n6308 ^ n6305;
  assign n6310 = ~n5962 & n6309;
  assign n6311 = n6310 ^ n6308;
  assign n6317 = x976 ^ x278;
  assign n6318 = n5970 & n6317;
  assign n6319 = n6318 ^ x278;
  assign n6312 = x1132 & n5989;
  assign n6313 = x1134 & n5986;
  assign n6314 = ~n6312 & ~n6313;
  assign n6315 = x1133 & n5993;
  assign n6316 = n6314 & ~n6315;
  assign n6320 = n6319 ^ n6316;
  assign n6321 = ~n5962 & ~n6320;
  assign n6322 = n6321 ^ n6319;
  assign n6328 = x958 ^ x279;
  assign n6329 = n5970 & n6328;
  assign n6330 = n6329 ^ x279;
  assign n6323 = x1133 & n5989;
  assign n6324 = x1135 & n5986;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = x1134 & n5993;
  assign n6327 = n6325 & ~n6326;
  assign n6331 = n6330 ^ n6327;
  assign n6332 = ~n5962 & ~n6331;
  assign n6333 = n6332 ^ n6330;
  assign n6339 = x914 ^ x280;
  assign n6340 = n5970 & ~n6339;
  assign n6341 = n6340 ^ x280;
  assign n6334 = x1135 & n5989;
  assign n6335 = x1137 & n5986;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = x1136 & n5993;
  assign n6338 = n6336 & ~n6337;
  assign n6342 = n6341 ^ n6338;
  assign n6343 = ~n5962 & n6342;
  assign n6344 = n6343 ^ n6341;
  assign n6350 = x830 ^ x281;
  assign n6351 = n5970 & ~n6350;
  assign n6352 = n6351 ^ x281;
  assign n6345 = x1137 & n5989;
  assign n6346 = x1139 & n5986;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = x1138 & n5993;
  assign n6349 = n6347 & ~n6348;
  assign n6353 = n6352 ^ n6349;
  assign n6354 = ~n5962 & n6353;
  assign n6355 = n6354 ^ n6352;
  assign n6361 = x836 ^ x282;
  assign n6362 = n5970 & ~n6361;
  assign n6363 = n6362 ^ x282;
  assign n6356 = x1138 & n5989;
  assign n6357 = x1140 & n5986;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = x1139 & n5993;
  assign n6360 = n6358 & ~n6359;
  assign n6364 = n6363 ^ n6360;
  assign n6365 = ~n5962 & n6364;
  assign n6366 = n6365 ^ n6363;
  assign n6368 = x1149 & n5986;
  assign n6369 = x1147 & n5989;
  assign n6370 = ~n6368 & ~n6369;
  assign n6371 = x1148 & n5993;
  assign n6372 = n6370 & ~n6371;
  assign n6367 = n5974 ^ x283;
  assign n6373 = n6372 ^ n6367;
  assign n6374 = ~n5962 & ~n6373;
  assign n6375 = n6374 ^ n6367;
  assign n6376 = x1143 & ~n3486;
  assign n6377 = n6376 ^ x284;
  assign n6378 = n6377 ^ x284;
  assign n6379 = n5685 ^ x284;
  assign n6380 = n6379 ^ x284;
  assign n6381 = n6378 & n6380;
  assign n6382 = n6381 ^ x284;
  assign n6383 = ~n6154 & ~n6382;
  assign n6384 = n6383 ^ x284;
  assign n6385 = n3332 & n3459;
  assign n6386 = ~n2894 & n6385;
  assign n6387 = x289 & n6386;
  assign n6388 = x286 & x288;
  assign n6389 = n6387 & n6388;
  assign n6390 = n6389 ^ x285;
  assign n6391 = ~x288 & n2894;
  assign n6392 = ~n6385 & n6391;
  assign n6393 = x285 & n2863;
  assign n6394 = n6392 & n6393;
  assign n6395 = ~x793 & ~n6394;
  assign n6396 = n6390 & n6395;
  assign n6397 = x288 & n6386;
  assign n6398 = n6397 ^ x286;
  assign n6399 = n6398 ^ n6392;
  assign n6400 = n2865 & ~n6398;
  assign n6401 = n6400 ^ x793;
  assign n6402 = ~n6399 & ~n6401;
  assign n6403 = n6402 ^ n6400;
  assign n6404 = ~x793 & n6403;
  assign n6405 = n6404 ^ x793;
  assign n6406 = ~x287 & x457;
  assign n6407 = ~x332 & ~n6406;
  assign n6408 = n2901 ^ x288;
  assign n6409 = n6408 ^ n6385;
  assign n6410 = ~x793 & n6409;
  assign n6411 = n6386 ^ x289;
  assign n6412 = n6411 ^ n6386;
  assign n6413 = n6397 ^ n6386;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = n6414 ^ n6386;
  assign n6416 = x286 & ~n6415;
  assign n6417 = x289 & ~n6388;
  assign n6418 = n6417 ^ n6393;
  assign n6419 = ~n6392 & n6418;
  assign n6420 = n6419 ^ n6393;
  assign n6421 = ~n6416 & ~n6420;
  assign n6422 = ~x793 & ~n6421;
  assign n6423 = x1048 ^ x290;
  assign n6424 = ~x476 & n6423;
  assign n6425 = n6424 ^ x290;
  assign n6426 = x1049 ^ x291;
  assign n6427 = ~x476 & n6426;
  assign n6428 = n6427 ^ x291;
  assign n6429 = x1084 ^ x292;
  assign n6430 = ~x476 & n6429;
  assign n6431 = n6430 ^ x292;
  assign n6432 = x1059 ^ x293;
  assign n6433 = ~x476 & n6432;
  assign n6434 = n6433 ^ x293;
  assign n6435 = x1072 ^ x294;
  assign n6436 = ~x476 & n6435;
  assign n6437 = n6436 ^ x294;
  assign n6438 = x1053 ^ x295;
  assign n6439 = ~x476 & n6438;
  assign n6440 = n6439 ^ x295;
  assign n6441 = x1037 ^ x296;
  assign n6442 = ~x476 & n6441;
  assign n6443 = n6442 ^ x296;
  assign n6444 = x1044 ^ x297;
  assign n6445 = ~x476 & n6444;
  assign n6446 = n6445 ^ x297;
  assign n6447 = x1044 ^ x298;
  assign n6448 = ~x478 & n6447;
  assign n6449 = n6448 ^ x298;
  assign n6450 = x106 & n3265;
  assign n6451 = x39 & ~x287;
  assign n6452 = n3490 & n6451;
  assign n6453 = ~n3495 & ~n6452;
  assign n6454 = ~n6450 & n6453;
  assign n6455 = n1571 & n1601;
  assign n6456 = n6454 & ~n6455;
  assign n6457 = ~x24 & n1579;
  assign n6458 = ~x312 & n6457;
  assign n6459 = n6458 ^ x300;
  assign n6460 = ~x55 & ~n6459;
  assign n6461 = ~x300 & ~x312;
  assign n6462 = n6457 & n6461;
  assign n6463 = n6462 ^ x301;
  assign n6464 = ~x55 & ~n6463;
  assign n6465 = n1776 ^ n1738;
  assign n6466 = n1729 & n6465;
  assign n6467 = n6466 ^ n1738;
  assign n6468 = x937 & n6467;
  assign n6469 = ~n1751 & ~n2215;
  assign n6470 = ~x237 & ~n6469;
  assign n6471 = ~n6468 & ~n6470;
  assign n6472 = n1779 ^ n1741;
  assign n6473 = n1729 & n6472;
  assign n6474 = n6473 ^ n1741;
  assign n6475 = x273 & n6474;
  assign n6476 = x1148 & ~n2294;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = n6471 & n6477;
  assign n6479 = x1049 ^ x303;
  assign n6480 = ~x478 & n6479;
  assign n6481 = n6480 ^ x303;
  assign n6482 = x1048 ^ x304;
  assign n6483 = ~x478 & n6482;
  assign n6484 = n6483 ^ x304;
  assign n6485 = x1084 ^ x305;
  assign n6486 = ~x478 & n6485;
  assign n6487 = n6486 ^ x305;
  assign n6488 = x1059 ^ x306;
  assign n6489 = ~x478 & n6488;
  assign n6490 = n6489 ^ x306;
  assign n6491 = x1053 ^ x307;
  assign n6492 = ~x478 & n6491;
  assign n6493 = n6492 ^ x307;
  assign n6494 = x1037 ^ x308;
  assign n6495 = ~x478 & n6494;
  assign n6496 = n6495 ^ x308;
  assign n6497 = x1072 ^ x309;
  assign n6498 = ~x478 & n6497;
  assign n6499 = n6498 ^ x309;
  assign n6500 = x271 & n6474;
  assign n6501 = ~x233 & ~n6469;
  assign n6502 = ~n6500 & ~n6501;
  assign n6503 = x1147 & ~n2294;
  assign n6504 = x934 & n6467;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = n6502 & n6505;
  assign n6507 = x301 & n6461;
  assign n6508 = n6457 & n6507;
  assign n6509 = n6508 ^ x311;
  assign n6510 = ~x55 & ~n6509;
  assign n6511 = n6457 ^ x312;
  assign n6512 = ~x55 & n6511;
  assign n6513 = n3921 ^ n2320;
  assign n6514 = n3921 ^ x314;
  assign n6515 = n6514 ^ x314;
  assign n6516 = n3908 ^ x314;
  assign n6517 = ~n6515 & n6516;
  assign n6518 = n6517 ^ x314;
  assign n6519 = n6513 & ~n6518;
  assign n6520 = n6519 ^ n2320;
  assign n6521 = n6520 ^ x313;
  assign n6522 = ~x954 & ~n6521;
  assign n6523 = n6522 ^ x313;
  assign n6524 = n4107 & n4414;
  assign n6525 = n4336 & n6524;
  assign n6526 = ~x340 & n6385;
  assign n6527 = x1080 ^ x315;
  assign n6528 = n6526 & n6527;
  assign n6529 = n6528 ^ x315;
  assign n6530 = x1047 ^ x316;
  assign n6531 = n6526 & n6530;
  assign n6532 = n6531 ^ x316;
  assign n6533 = ~x330 & n6385;
  assign n6534 = x1078 ^ x317;
  assign n6535 = n6533 & n6534;
  assign n6536 = n6535 ^ x317;
  assign n6537 = ~x341 & n6385;
  assign n6538 = x1074 ^ x318;
  assign n6539 = n6537 & n6538;
  assign n6540 = n6539 ^ x318;
  assign n6541 = x1072 ^ x319;
  assign n6542 = n6537 & n6541;
  assign n6543 = n6542 ^ x319;
  assign n6544 = x1048 ^ x320;
  assign n6545 = n6526 & n6544;
  assign n6546 = n6545 ^ x320;
  assign n6547 = x1058 ^ x321;
  assign n6548 = n6526 & n6547;
  assign n6549 = n6548 ^ x321;
  assign n6550 = x1051 ^ x322;
  assign n6551 = n6526 & n6550;
  assign n6552 = n6551 ^ x322;
  assign n6553 = x1065 ^ x323;
  assign n6554 = n6526 & n6553;
  assign n6555 = n6554 ^ x323;
  assign n6556 = x1086 ^ x324;
  assign n6557 = n6537 & n6556;
  assign n6558 = n6557 ^ x324;
  assign n6559 = x1063 ^ x325;
  assign n6560 = n6537 & n6559;
  assign n6561 = n6560 ^ x325;
  assign n6562 = x1057 ^ x326;
  assign n6563 = n6537 & n6562;
  assign n6564 = n6563 ^ x326;
  assign n6565 = x1040 ^ x327;
  assign n6566 = n6526 & n6565;
  assign n6567 = n6566 ^ x327;
  assign n6568 = x1058 ^ x328;
  assign n6569 = n6537 & n6568;
  assign n6570 = n6569 ^ x328;
  assign n6571 = x1043 ^ x329;
  assign n6572 = n6537 & n6571;
  assign n6573 = n6572 ^ x329;
  assign n6574 = x1092 & ~n1471;
  assign n6575 = x340 ^ x330;
  assign n6576 = n6385 & n6575;
  assign n6577 = n6576 ^ x330;
  assign n6578 = n6574 & ~n6577;
  assign n6579 = x341 ^ x331;
  assign n6580 = n6385 & n6579;
  assign n6581 = n6580 ^ x331;
  assign n6582 = n6574 & ~n6581;
  assign n6583 = n1752 & n3268;
  assign n6584 = ~n3424 & ~n3582;
  assign n6585 = ~n1588 & n6584;
  assign n6586 = ~n6583 & n6585;
  assign n6587 = x1040 ^ x333;
  assign n6588 = n6537 & n6587;
  assign n6589 = n6588 ^ x333;
  assign n6590 = x1065 ^ x334;
  assign n6591 = n6537 & n6590;
  assign n6592 = n6591 ^ x334;
  assign n6593 = x1069 ^ x335;
  assign n6594 = n6537 & n6593;
  assign n6595 = n6594 ^ x335;
  assign n6596 = x1070 ^ x336;
  assign n6597 = n6533 & n6596;
  assign n6598 = n6597 ^ x336;
  assign n6599 = x1044 ^ x337;
  assign n6600 = n6533 & n6599;
  assign n6601 = n6600 ^ x337;
  assign n6602 = x1072 ^ x338;
  assign n6603 = n6533 & n6602;
  assign n6604 = n6603 ^ x338;
  assign n6605 = x1086 ^ x339;
  assign n6606 = n6533 & n6605;
  assign n6607 = n6606 ^ x339;
  assign n6608 = n6385 ^ x340;
  assign n6609 = n6608 ^ x340;
  assign n6610 = x340 ^ x331;
  assign n6611 = n6609 & n6610;
  assign n6612 = n6611 ^ x340;
  assign n6613 = n6574 & n6612;
  assign n6614 = x341 ^ x330;
  assign n6615 = ~n6385 & n6614;
  assign n6616 = n6615 ^ x330;
  assign n6617 = n6574 & ~n6616;
  assign n6618 = x1049 ^ x342;
  assign n6619 = n6526 & n6618;
  assign n6620 = n6619 ^ x342;
  assign n6621 = x1062 ^ x343;
  assign n6622 = n6526 & n6621;
  assign n6623 = n6622 ^ x343;
  assign n6624 = x1069 ^ x344;
  assign n6625 = n6526 & n6624;
  assign n6626 = n6625 ^ x344;
  assign n6627 = x1039 ^ x345;
  assign n6628 = n6526 & n6627;
  assign n6629 = n6628 ^ x345;
  assign n6630 = x1067 ^ x346;
  assign n6631 = n6526 & n6630;
  assign n6632 = n6631 ^ x346;
  assign n6633 = x1055 ^ x347;
  assign n6634 = n6526 & n6633;
  assign n6635 = n6634 ^ x347;
  assign n6636 = x1087 ^ x348;
  assign n6637 = n6526 & n6636;
  assign n6638 = n6637 ^ x348;
  assign n6639 = x1043 ^ x349;
  assign n6640 = n6526 & n6639;
  assign n6641 = n6640 ^ x349;
  assign n6642 = x1035 ^ x350;
  assign n6643 = n6526 & n6642;
  assign n6644 = n6643 ^ x350;
  assign n6645 = x1079 ^ x351;
  assign n6646 = n6526 & n6645;
  assign n6647 = n6646 ^ x351;
  assign n6648 = x1078 ^ x352;
  assign n6649 = n6526 & n6648;
  assign n6650 = n6649 ^ x352;
  assign n6651 = x1063 ^ x353;
  assign n6652 = n6526 & n6651;
  assign n6653 = n6652 ^ x353;
  assign n6654 = x1045 ^ x354;
  assign n6655 = n6526 & n6654;
  assign n6656 = n6655 ^ x354;
  assign n6657 = x1084 ^ x355;
  assign n6658 = n6526 & n6657;
  assign n6659 = n6658 ^ x355;
  assign n6660 = x1081 ^ x356;
  assign n6661 = n6526 & n6660;
  assign n6662 = n6661 ^ x356;
  assign n6663 = x1076 ^ x357;
  assign n6664 = n6526 & n6663;
  assign n6665 = n6664 ^ x357;
  assign n6666 = x1071 ^ x358;
  assign n6667 = n6526 & n6666;
  assign n6668 = n6667 ^ x358;
  assign n6669 = x1068 ^ x359;
  assign n6670 = n6526 & n6669;
  assign n6671 = n6670 ^ x359;
  assign n6672 = x1042 ^ x360;
  assign n6673 = n6526 & n6672;
  assign n6674 = n6673 ^ x360;
  assign n6675 = x1059 ^ x361;
  assign n6676 = n6526 & n6675;
  assign n6677 = n6676 ^ x361;
  assign n6678 = x1070 ^ x362;
  assign n6679 = n6526 & n6678;
  assign n6680 = n6679 ^ x362;
  assign n6681 = x1049 ^ x363;
  assign n6682 = n6533 & n6681;
  assign n6683 = n6682 ^ x363;
  assign n6684 = x1062 ^ x364;
  assign n6685 = n6533 & n6684;
  assign n6686 = n6685 ^ x364;
  assign n6687 = x1065 ^ x365;
  assign n6688 = n6533 & n6687;
  assign n6689 = n6688 ^ x365;
  assign n6690 = x1069 ^ x366;
  assign n6691 = n6533 & n6690;
  assign n6692 = n6691 ^ x366;
  assign n6693 = x1039 ^ x367;
  assign n6694 = n6533 & n6693;
  assign n6695 = n6694 ^ x367;
  assign n6696 = x1067 ^ x368;
  assign n6697 = n6533 & n6696;
  assign n6698 = n6697 ^ x368;
  assign n6699 = x1080 ^ x369;
  assign n6700 = n6533 & n6699;
  assign n6701 = n6700 ^ x369;
  assign n6702 = x1055 ^ x370;
  assign n6703 = n6533 & n6702;
  assign n6704 = n6703 ^ x370;
  assign n6705 = x1051 ^ x371;
  assign n6706 = n6533 & n6705;
  assign n6707 = n6706 ^ x371;
  assign n6708 = x1048 ^ x372;
  assign n6709 = n6533 & n6708;
  assign n6710 = n6709 ^ x372;
  assign n6711 = x1087 ^ x373;
  assign n6712 = n6533 & n6711;
  assign n6713 = n6712 ^ x373;
  assign n6714 = x1035 ^ x374;
  assign n6715 = n6533 & n6714;
  assign n6716 = n6715 ^ x374;
  assign n6717 = x1047 ^ x375;
  assign n6718 = n6533 & n6717;
  assign n6719 = n6718 ^ x375;
  assign n6720 = x1079 ^ x376;
  assign n6721 = n6533 & n6720;
  assign n6722 = n6721 ^ x376;
  assign n6723 = x1074 ^ x377;
  assign n6724 = n6533 & n6723;
  assign n6725 = n6724 ^ x377;
  assign n6726 = x1063 ^ x378;
  assign n6727 = n6533 & n6726;
  assign n6728 = n6727 ^ x378;
  assign n6729 = x1045 ^ x379;
  assign n6730 = n6533 & n6729;
  assign n6731 = n6730 ^ x379;
  assign n6732 = x1084 ^ x380;
  assign n6733 = n6533 & n6732;
  assign n6734 = n6733 ^ x380;
  assign n6735 = x1081 ^ x381;
  assign n6736 = n6533 & n6735;
  assign n6737 = n6736 ^ x381;
  assign n6738 = x1076 ^ x382;
  assign n6739 = n6533 & n6738;
  assign n6740 = n6739 ^ x382;
  assign n6741 = x1071 ^ x383;
  assign n6742 = n6533 & n6741;
  assign n6743 = n6742 ^ x383;
  assign n6744 = x1068 ^ x384;
  assign n6745 = n6533 & n6744;
  assign n6746 = n6745 ^ x384;
  assign n6747 = x1042 ^ x385;
  assign n6748 = n6533 & n6747;
  assign n6749 = n6748 ^ x385;
  assign n6750 = x1059 ^ x386;
  assign n6751 = n6533 & n6750;
  assign n6752 = n6751 ^ x386;
  assign n6753 = x1053 ^ x387;
  assign n6754 = n6533 & n6753;
  assign n6755 = n6754 ^ x387;
  assign n6756 = x1037 ^ x388;
  assign n6757 = n6533 & n6756;
  assign n6758 = n6757 ^ x388;
  assign n6759 = x1036 ^ x389;
  assign n6760 = n6533 & n6759;
  assign n6761 = n6760 ^ x389;
  assign n6762 = x1049 ^ x390;
  assign n6763 = n6537 & n6762;
  assign n6764 = n6763 ^ x390;
  assign n6765 = x1062 ^ x391;
  assign n6766 = n6537 & n6765;
  assign n6767 = n6766 ^ x391;
  assign n6768 = x1039 ^ x392;
  assign n6769 = n6537 & n6768;
  assign n6770 = n6769 ^ x392;
  assign n6771 = x1067 ^ x393;
  assign n6772 = n6537 & n6771;
  assign n6773 = n6772 ^ x393;
  assign n6774 = x1080 ^ x394;
  assign n6775 = n6537 & n6774;
  assign n6776 = n6775 ^ x394;
  assign n6777 = x1055 ^ x395;
  assign n6778 = n6537 & n6777;
  assign n6779 = n6778 ^ x395;
  assign n6780 = x1051 ^ x396;
  assign n6781 = n6537 & n6780;
  assign n6782 = n6781 ^ x396;
  assign n6783 = x1048 ^ x397;
  assign n6784 = n6537 & n6783;
  assign n6785 = n6784 ^ x397;
  assign n6786 = x1087 ^ x398;
  assign n6787 = n6537 & n6786;
  assign n6788 = n6787 ^ x398;
  assign n6789 = x1047 ^ x399;
  assign n6790 = n6537 & n6789;
  assign n6791 = n6790 ^ x399;
  assign n6792 = x1035 ^ x400;
  assign n6793 = n6537 & n6792;
  assign n6794 = n6793 ^ x400;
  assign n6795 = x1079 ^ x401;
  assign n6796 = n6537 & n6795;
  assign n6797 = n6796 ^ x401;
  assign n6798 = x1078 ^ x402;
  assign n6799 = n6537 & n6798;
  assign n6800 = n6799 ^ x402;
  assign n6801 = x1045 ^ x403;
  assign n6802 = n6537 & n6801;
  assign n6803 = n6802 ^ x403;
  assign n6804 = x1084 ^ x404;
  assign n6805 = n6537 & n6804;
  assign n6806 = n6805 ^ x404;
  assign n6807 = x1081 ^ x405;
  assign n6808 = n6537 & n6807;
  assign n6809 = n6808 ^ x405;
  assign n6810 = x1076 ^ x406;
  assign n6811 = n6537 & n6810;
  assign n6812 = n6811 ^ x406;
  assign n6813 = x1071 ^ x407;
  assign n6814 = n6537 & n6813;
  assign n6815 = n6814 ^ x407;
  assign n6816 = x1068 ^ x408;
  assign n6817 = n6537 & n6816;
  assign n6818 = n6817 ^ x408;
  assign n6819 = x1042 ^ x409;
  assign n6820 = n6537 & n6819;
  assign n6821 = n6820 ^ x409;
  assign n6822 = x1059 ^ x410;
  assign n6823 = n6537 & n6822;
  assign n6824 = n6823 ^ x410;
  assign n6825 = x1053 ^ x411;
  assign n6826 = n6537 & n6825;
  assign n6827 = n6826 ^ x411;
  assign n6828 = x1037 ^ x412;
  assign n6829 = n6537 & n6828;
  assign n6830 = n6829 ^ x412;
  assign n6831 = x1036 ^ x413;
  assign n6832 = n6537 & n6831;
  assign n6833 = n6832 ^ x413;
  assign n6834 = ~x331 & n6385;
  assign n6835 = x1049 ^ x414;
  assign n6836 = n6834 & n6835;
  assign n6837 = n6836 ^ x414;
  assign n6838 = x1062 ^ x415;
  assign n6839 = n6834 & n6838;
  assign n6840 = n6839 ^ x415;
  assign n6841 = x1069 ^ x416;
  assign n6842 = n6834 & n6841;
  assign n6843 = n6842 ^ x416;
  assign n6844 = x1039 ^ x417;
  assign n6845 = n6834 & n6844;
  assign n6846 = n6845 ^ x417;
  assign n6847 = x1067 ^ x418;
  assign n6848 = n6834 & n6847;
  assign n6849 = n6848 ^ x418;
  assign n6850 = x1080 ^ x419;
  assign n6851 = n6834 & n6850;
  assign n6852 = n6851 ^ x419;
  assign n6853 = x1055 ^ x420;
  assign n6854 = n6834 & n6853;
  assign n6855 = n6854 ^ x420;
  assign n6856 = x1051 ^ x421;
  assign n6857 = n6834 & n6856;
  assign n6858 = n6857 ^ x421;
  assign n6859 = x1048 ^ x422;
  assign n6860 = n6834 & n6859;
  assign n6861 = n6860 ^ x422;
  assign n6862 = x1087 ^ x423;
  assign n6863 = n6834 & n6862;
  assign n6864 = n6863 ^ x423;
  assign n6865 = x1047 ^ x424;
  assign n6866 = n6834 & n6865;
  assign n6867 = n6866 ^ x424;
  assign n6868 = x1035 ^ x425;
  assign n6869 = n6834 & n6868;
  assign n6870 = n6869 ^ x425;
  assign n6871 = x1079 ^ x426;
  assign n6872 = n6834 & n6871;
  assign n6873 = n6872 ^ x426;
  assign n6874 = x1078 ^ x427;
  assign n6875 = n6834 & n6874;
  assign n6876 = n6875 ^ x427;
  assign n6877 = x1045 ^ x428;
  assign n6878 = n6834 & n6877;
  assign n6879 = n6878 ^ x428;
  assign n6880 = x1084 ^ x429;
  assign n6881 = n6834 & n6880;
  assign n6882 = n6881 ^ x429;
  assign n6883 = x1076 ^ x430;
  assign n6884 = n6834 & n6883;
  assign n6885 = n6884 ^ x430;
  assign n6886 = x1071 ^ x431;
  assign n6887 = n6834 & n6886;
  assign n6888 = n6887 ^ x431;
  assign n6889 = x1068 ^ x432;
  assign n6890 = n6834 & n6889;
  assign n6891 = n6890 ^ x432;
  assign n6892 = x1042 ^ x433;
  assign n6893 = n6834 & n6892;
  assign n6894 = n6893 ^ x433;
  assign n6895 = x1059 ^ x434;
  assign n6896 = n6834 & n6895;
  assign n6897 = n6896 ^ x434;
  assign n6898 = x1053 ^ x435;
  assign n6899 = n6834 & n6898;
  assign n6900 = n6899 ^ x435;
  assign n6901 = x1037 ^ x436;
  assign n6902 = n6834 & n6901;
  assign n6903 = n6902 ^ x436;
  assign n6904 = x1070 ^ x437;
  assign n6905 = n6834 & n6904;
  assign n6906 = n6905 ^ x437;
  assign n6907 = x1036 ^ x438;
  assign n6908 = n6834 & n6907;
  assign n6909 = n6908 ^ x438;
  assign n6910 = x1057 ^ x439;
  assign n6911 = n6533 & n6910;
  assign n6912 = n6911 ^ x439;
  assign n6913 = x1043 ^ x440;
  assign n6914 = n6533 & n6913;
  assign n6915 = n6914 ^ x440;
  assign n6916 = x1044 ^ x441;
  assign n6917 = n6526 & n6916;
  assign n6918 = n6917 ^ x441;
  assign n6919 = x1058 ^ x442;
  assign n6920 = n6533 & n6919;
  assign n6921 = n6920 ^ x442;
  assign n6922 = x1044 ^ x443;
  assign n6923 = n6834 & n6922;
  assign n6924 = n6923 ^ x443;
  assign n6925 = x1072 ^ x444;
  assign n6926 = n6834 & n6925;
  assign n6927 = n6926 ^ x444;
  assign n6928 = x1081 ^ x445;
  assign n6929 = n6834 & n6928;
  assign n6930 = n6929 ^ x445;
  assign n6931 = x1086 ^ x446;
  assign n6932 = n6834 & n6931;
  assign n6933 = n6932 ^ x446;
  assign n6934 = x1040 ^ x447;
  assign n6935 = n6533 & n6934;
  assign n6936 = n6935 ^ x447;
  assign n6937 = x1074 ^ x448;
  assign n6938 = n6834 & n6937;
  assign n6939 = n6938 ^ x448;
  assign n6940 = x1057 ^ x449;
  assign n6941 = n6834 & n6940;
  assign n6942 = n6941 ^ x449;
  assign n6943 = x1036 ^ x450;
  assign n6944 = n6526 & n6943;
  assign n6945 = n6944 ^ x450;
  assign n6946 = x1063 ^ x451;
  assign n6947 = n6834 & n6946;
  assign n6948 = n6947 ^ x451;
  assign n6949 = x1053 ^ x452;
  assign n6950 = n6526 & n6949;
  assign n6951 = n6950 ^ x452;
  assign n6952 = x1040 ^ x453;
  assign n6953 = n6834 & n6952;
  assign n6954 = n6953 ^ x453;
  assign n6955 = x1043 ^ x454;
  assign n6956 = n6834 & n6955;
  assign n6957 = n6956 ^ x454;
  assign n6958 = x1037 ^ x455;
  assign n6959 = n6526 & n6958;
  assign n6960 = n6959 ^ x455;
  assign n6961 = x1044 ^ x456;
  assign n6962 = n6537 & n6961;
  assign n6963 = n6962 ^ x456;
  assign n6964 = x599 & x815;
  assign n6965 = x810 & ~n6964;
  assign n6966 = x596 & ~n6965;
  assign n6967 = x804 & ~n6966;
  assign n6968 = x594 & x600;
  assign n6969 = x597 & x601;
  assign n6970 = n6968 & n6969;
  assign n6971 = ~x804 & ~x810;
  assign n6972 = ~x595 & ~n6971;
  assign n6973 = n6970 & ~n6972;
  assign n6974 = ~n6967 & n6973;
  assign n6975 = ~x601 & ~n6971;
  assign n6976 = ~x815 & ~n6975;
  assign n6977 = x600 & ~x810;
  assign n6978 = x804 & ~n6977;
  assign n6979 = n6976 & ~n6978;
  assign n6980 = ~n6974 & ~n6979;
  assign n6981 = x605 & ~n6980;
  assign n6982 = ~x815 & x990;
  assign n6983 = n6968 & n6982;
  assign n6984 = n6978 & n6983;
  assign n6985 = ~n6981 & ~n6984;
  assign n6986 = x821 & ~n6985;
  assign n6987 = x1072 ^ x458;
  assign n6988 = n6526 & n6987;
  assign n6989 = n6988 ^ x458;
  assign n6990 = x1058 ^ x459;
  assign n6991 = n6834 & n6990;
  assign n6992 = n6991 ^ x459;
  assign n6993 = x1086 ^ x460;
  assign n6994 = n6526 & n6993;
  assign n6995 = n6994 ^ x460;
  assign n6996 = x1057 ^ x461;
  assign n6997 = n6526 & n6996;
  assign n6998 = n6997 ^ x461;
  assign n6999 = x1074 ^ x462;
  assign n7000 = n6526 & n6999;
  assign n7001 = n7000 ^ x462;
  assign n7002 = x1070 ^ x463;
  assign n7003 = n6537 & n7002;
  assign n7004 = n7003 ^ x463;
  assign n7005 = x1065 ^ x464;
  assign n7006 = n6834 & n7005;
  assign n7007 = n7006 ^ x464;
  assign n7008 = ~x243 & n6474;
  assign n7009 = x926 & n6467;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = x1157 & ~n2294;
  assign n7012 = n7010 & ~n7011;
  assign n7013 = x275 & n6474;
  assign n7014 = x943 & n6467;
  assign n7015 = ~n7013 & ~n7014;
  assign n7016 = x1151 & ~n2294;
  assign n7017 = n7015 & ~n7016;
  assign n7018 = n3547 & n5526;
  assign n7019 = x40 & x1001;
  assign n7020 = n2381 & n7019;
  assign n7021 = n2390 & n7020;
  assign n7022 = ~n7018 & ~n7021;
  assign n7023 = ~x24 & n1588;
  assign n7024 = x468 & ~n7023;
  assign n7025 = ~n3525 & ~n7024;
  assign n7026 = x942 & n6467;
  assign n7027 = ~x263 & n6474;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = x1156 & ~n2294;
  assign n7030 = n7028 & ~n7029;
  assign n7031 = x925 & n6467;
  assign n7032 = x267 & n6474;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = x1155 & ~n2294;
  assign n7035 = n7033 & ~n7034;
  assign n7036 = x941 & n6467;
  assign n7037 = x253 & n6474;
  assign n7038 = ~n7036 & ~n7037;
  assign n7039 = x1153 & ~n2294;
  assign n7040 = n7038 & ~n7039;
  assign n7041 = x254 & n6474;
  assign n7042 = x923 & n6467;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = x1154 & ~n2294;
  assign n7045 = n7043 & ~n7044;
  assign n7046 = x922 & n6467;
  assign n7047 = x268 & n6474;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = x1152 & ~n2294;
  assign n7050 = n7048 & ~n7049;
  assign n7051 = x931 & n6467;
  assign n7052 = x272 & n6474;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = x1150 & ~n2294;
  assign n7055 = n7053 & ~n7054;
  assign n7056 = x936 & n6467;
  assign n7057 = x283 & n6474;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = x1149 & ~n2294;
  assign n7060 = n7058 & ~n7059;
  assign n7061 = x71 & n5993;
  assign n7062 = ~n3788 & ~n7061;
  assign n7063 = x71 & n5989;
  assign n7064 = x481 ^ x248;
  assign n7065 = ~n5274 & n7064;
  assign n7066 = n7065 ^ x248;
  assign n7067 = x482 ^ x249;
  assign n7068 = ~n5289 & n7067;
  assign n7069 = n7068 ^ x249;
  assign n7070 = x483 ^ x242;
  assign n7071 = ~n5314 & n7070;
  assign n7072 = n7071 ^ x242;
  assign n7073 = x484 ^ x249;
  assign n7074 = ~n5314 & n7073;
  assign n7075 = n7074 ^ x249;
  assign n7076 = x485 ^ x234;
  assign n7077 = ~n5429 & n7076;
  assign n7078 = n7077 ^ x234;
  assign n7079 = x486 ^ x244;
  assign n7080 = ~n5429 & n7079;
  assign n7081 = n7080 ^ x244;
  assign n7082 = x487 ^ x246;
  assign n7083 = ~n5274 & n7082;
  assign n7084 = n7083 ^ x246;
  assign n7085 = x488 ^ x239;
  assign n7086 = ~n5274 & ~n7085;
  assign n7087 = n7086 ^ x239;
  assign n7088 = x489 ^ x242;
  assign n7089 = ~n5429 & n7088;
  assign n7090 = n7089 ^ x242;
  assign n7091 = x490 ^ x241;
  assign n7092 = ~n5314 & n7091;
  assign n7093 = n7092 ^ x241;
  assign n7094 = x491 ^ x238;
  assign n7095 = ~n5314 & n7094;
  assign n7096 = n7095 ^ x238;
  assign n7097 = x492 ^ x240;
  assign n7098 = ~n5314 & n7097;
  assign n7099 = n7098 ^ x240;
  assign n7100 = x493 ^ x244;
  assign n7101 = ~n5314 & n7100;
  assign n7102 = n7101 ^ x244;
  assign n7103 = x494 ^ x239;
  assign n7104 = ~n5314 & ~n7103;
  assign n7105 = n7104 ^ x239;
  assign n7106 = x495 ^ x235;
  assign n7107 = ~n5314 & n7106;
  assign n7108 = n7107 ^ x235;
  assign n7109 = x496 ^ x249;
  assign n7110 = ~n5307 & n7109;
  assign n7111 = n7110 ^ x249;
  assign n7112 = x497 ^ x239;
  assign n7113 = ~n5307 & ~n7112;
  assign n7114 = n7113 ^ x239;
  assign n7115 = x498 ^ x238;
  assign n7116 = ~n5289 & n7115;
  assign n7117 = n7116 ^ x238;
  assign n7118 = x499 ^ x246;
  assign n7119 = ~n5307 & n7118;
  assign n7120 = n7119 ^ x246;
  assign n7121 = x500 ^ x241;
  assign n7122 = ~n5307 & n7121;
  assign n7123 = n7122 ^ x241;
  assign n7124 = x501 ^ x248;
  assign n7125 = ~n5307 & n7124;
  assign n7126 = n7125 ^ x248;
  assign n7127 = x502 ^ x247;
  assign n7128 = ~n5307 & n7127;
  assign n7129 = n7128 ^ x247;
  assign n7130 = x503 ^ x245;
  assign n7131 = ~n5307 & n7130;
  assign n7132 = n7131 ^ x245;
  assign n7133 = x504 ^ x242;
  assign n7134 = ~n5303 & n7133;
  assign n7135 = n7134 ^ x242;
  assign n7136 = x505 ^ x234;
  assign n7137 = ~n5307 & n7136;
  assign n7138 = n7137 ^ x234;
  assign n7139 = x506 ^ x241;
  assign n7140 = ~n5303 & n7139;
  assign n7141 = n7140 ^ x241;
  assign n7142 = x507 ^ x238;
  assign n7143 = ~n5303 & n7142;
  assign n7144 = n7143 ^ x238;
  assign n7145 = x508 ^ x247;
  assign n7146 = ~n5303 & n7145;
  assign n7147 = n7146 ^ x247;
  assign n7148 = x509 ^ x245;
  assign n7149 = ~n5303 & n7148;
  assign n7150 = n7149 ^ x245;
  assign n7151 = x510 ^ x242;
  assign n7152 = ~n5274 & n7151;
  assign n7153 = n7152 ^ x242;
  assign n7154 = x511 ^ x234;
  assign n7155 = ~n5274 & n7154;
  assign n7156 = n7155 ^ x234;
  assign n7157 = x512 ^ x235;
  assign n7158 = ~n5274 & n7157;
  assign n7159 = n7158 ^ x235;
  assign n7160 = x513 ^ x244;
  assign n7161 = ~n5274 & n7160;
  assign n7162 = n7161 ^ x244;
  assign n7163 = x514 ^ x245;
  assign n7164 = ~n5274 & n7163;
  assign n7165 = n7164 ^ x245;
  assign n7166 = x515 ^ x240;
  assign n7167 = ~n5274 & n7166;
  assign n7168 = n7167 ^ x240;
  assign n7169 = x516 ^ x247;
  assign n7170 = ~n5274 & n7169;
  assign n7171 = n7170 ^ x247;
  assign n7172 = x517 ^ x238;
  assign n7173 = ~n5274 & n7172;
  assign n7174 = n7173 ^ x238;
  assign n7175 = x518 ^ x234;
  assign n7176 = ~n5282 & n7175;
  assign n7177 = n7176 ^ x234;
  assign n7178 = x519 ^ x239;
  assign n7179 = ~n5282 & ~n7178;
  assign n7180 = n7179 ^ x239;
  assign n7181 = x520 ^ x246;
  assign n7182 = ~n5282 & n7181;
  assign n7183 = n7182 ^ x246;
  assign n7184 = x521 ^ x248;
  assign n7185 = ~n5282 & n7184;
  assign n7186 = n7185 ^ x248;
  assign n7187 = x522 ^ x238;
  assign n7188 = ~n5282 & n7187;
  assign n7189 = n7188 ^ x238;
  assign n7190 = x523 ^ x234;
  assign n7191 = ~n5442 & n7190;
  assign n7192 = n7191 ^ x234;
  assign n7193 = x524 ^ x239;
  assign n7194 = ~n5442 & ~n7193;
  assign n7195 = n7194 ^ x239;
  assign n7196 = x525 ^ x245;
  assign n7197 = ~n5442 & n7196;
  assign n7198 = n7197 ^ x245;
  assign n7199 = x526 ^ x246;
  assign n7200 = ~n5442 & n7199;
  assign n7201 = n7200 ^ x246;
  assign n7202 = x527 ^ x247;
  assign n7203 = ~n5442 & n7202;
  assign n7204 = n7203 ^ x247;
  assign n7205 = x528 ^ x249;
  assign n7206 = ~n5442 & n7205;
  assign n7207 = n7206 ^ x249;
  assign n7208 = x529 ^ x238;
  assign n7209 = ~n5442 & n7208;
  assign n7210 = n7209 ^ x238;
  assign n7211 = x530 ^ x240;
  assign n7212 = ~n5442 & n7211;
  assign n7213 = n7212 ^ x240;
  assign n7214 = x531 ^ x235;
  assign n7215 = ~n5289 & n7214;
  assign n7216 = n7215 ^ x235;
  assign n7217 = x532 ^ x247;
  assign n7218 = ~n5289 & n7217;
  assign n7219 = n7218 ^ x247;
  assign n7220 = x533 ^ x235;
  assign n7221 = ~n5303 & n7220;
  assign n7222 = n7221 ^ x235;
  assign n7223 = x534 ^ x239;
  assign n7224 = ~n5303 & ~n7223;
  assign n7225 = n7224 ^ x239;
  assign n7226 = x535 ^ x240;
  assign n7227 = ~n5303 & n7226;
  assign n7228 = n7227 ^ x240;
  assign n7229 = x536 ^ x246;
  assign n7230 = ~n5303 & n7229;
  assign n7231 = n7230 ^ x246;
  assign n7232 = x537 ^ x248;
  assign n7233 = ~n5303 & n7232;
  assign n7234 = n7233 ^ x248;
  assign n7235 = x538 ^ x249;
  assign n7236 = ~n5303 & n7235;
  assign n7237 = n7236 ^ x249;
  assign n7238 = x539 ^ x242;
  assign n7239 = ~n5307 & n7238;
  assign n7240 = n7239 ^ x242;
  assign n7241 = x540 ^ x235;
  assign n7242 = ~n5307 & n7241;
  assign n7243 = n7242 ^ x235;
  assign n7244 = x541 ^ x244;
  assign n7245 = ~n5307 & n7244;
  assign n7246 = n7245 ^ x244;
  assign n7247 = x542 ^ x240;
  assign n7248 = ~n5307 & n7247;
  assign n7249 = n7248 ^ x240;
  assign n7250 = x543 ^ x238;
  assign n7251 = ~n5307 & n7250;
  assign n7252 = n7251 ^ x238;
  assign n7253 = x544 ^ x234;
  assign n7254 = ~n5314 & n7253;
  assign n7255 = n7254 ^ x234;
  assign n7256 = x545 ^ x245;
  assign n7257 = ~n5314 & n7256;
  assign n7258 = n7257 ^ x245;
  assign n7259 = x546 ^ x246;
  assign n7260 = ~n5314 & n7259;
  assign n7261 = n7260 ^ x246;
  assign n7262 = x547 ^ x247;
  assign n7263 = ~n5314 & n7262;
  assign n7264 = n7263 ^ x247;
  assign n7265 = x548 ^ x248;
  assign n7266 = ~n5314 & n7265;
  assign n7267 = n7266 ^ x248;
  assign n7268 = x549 ^ x235;
  assign n7269 = ~n5429 & n7268;
  assign n7270 = n7269 ^ x235;
  assign n7271 = x550 ^ x239;
  assign n7272 = ~n5429 & ~n7271;
  assign n7273 = n7272 ^ x239;
  assign n7274 = x551 ^ x240;
  assign n7275 = ~n5429 & n7274;
  assign n7276 = n7275 ^ x240;
  assign n7277 = x552 ^ x247;
  assign n7278 = ~n5429 & n7277;
  assign n7279 = n7278 ^ x247;
  assign n7280 = x553 ^ x241;
  assign n7281 = ~n5429 & n7280;
  assign n7282 = n7281 ^ x241;
  assign n7283 = x554 ^ x248;
  assign n7284 = ~n5429 & n7283;
  assign n7285 = n7284 ^ x248;
  assign n7286 = x555 ^ x249;
  assign n7287 = ~n5429 & n7286;
  assign n7288 = n7287 ^ x249;
  assign n7289 = x556 ^ x242;
  assign n7290 = ~n5289 & n7289;
  assign n7291 = n7290 ^ x242;
  assign n7292 = x557 ^ x234;
  assign n7293 = ~n5303 & n7292;
  assign n7294 = n7293 ^ x234;
  assign n7295 = x558 ^ x244;
  assign n7296 = ~n5303 & n7295;
  assign n7297 = n7296 ^ x244;
  assign n7298 = x559 ^ x241;
  assign n7299 = ~n5274 & n7298;
  assign n7300 = n7299 ^ x241;
  assign n7301 = x560 ^ x240;
  assign n7302 = ~n5289 & n7301;
  assign n7303 = n7302 ^ x240;
  assign n7304 = x561 ^ x247;
  assign n7305 = ~n5282 & n7304;
  assign n7306 = n7305 ^ x247;
  assign n7307 = x562 ^ x241;
  assign n7308 = ~n5289 & n7307;
  assign n7309 = n7308 ^ x241;
  assign n7310 = x563 ^ x246;
  assign n7311 = ~n5429 & n7310;
  assign n7312 = n7311 ^ x246;
  assign n7313 = x564 ^ x246;
  assign n7314 = ~n5289 & n7313;
  assign n7315 = n7314 ^ x246;
  assign n7316 = x565 ^ x248;
  assign n7317 = ~n5289 & n7316;
  assign n7318 = n7317 ^ x248;
  assign n7319 = x566 ^ x244;
  assign n7320 = ~n5289 & n7319;
  assign n7321 = n7320 ^ x244;
  assign n7322 = x230 & x1093;
  assign n7323 = x1091 ^ x567;
  assign n7324 = n7323 ^ x567;
  assign n7325 = x665 & n4604;
  assign n7326 = x621 & n4578;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = n7327 ^ x567;
  assign n7329 = n7328 ^ x567;
  assign n7330 = n7324 & ~n7329;
  assign n7331 = n7330 ^ x567;
  assign n7332 = n7322 & ~n7331;
  assign n7333 = n7332 ^ x567;
  assign n7334 = x1092 & ~n7333;
  assign n7335 = x568 ^ x245;
  assign n7336 = ~n5289 & n7335;
  assign n7337 = n7336 ^ x245;
  assign n7338 = x569 ^ x239;
  assign n7339 = ~n5289 & ~n7338;
  assign n7340 = n7339 ^ x239;
  assign n7341 = x570 ^ x234;
  assign n7342 = ~n5289 & n7341;
  assign n7343 = n7342 ^ x234;
  assign n7344 = x571 ^ x241;
  assign n7345 = ~n5442 & n7344;
  assign n7346 = n7345 ^ x241;
  assign n7347 = x572 ^ x244;
  assign n7348 = ~n5442 & n7347;
  assign n7349 = n7348 ^ x244;
  assign n7350 = x573 ^ x242;
  assign n7351 = ~n5442 & n7350;
  assign n7352 = n7351 ^ x242;
  assign n7353 = x574 ^ x241;
  assign n7354 = ~n5282 & n7353;
  assign n7355 = n7354 ^ x241;
  assign n7356 = x575 ^ x235;
  assign n7357 = ~n5442 & n7356;
  assign n7358 = n7357 ^ x235;
  assign n7359 = x576 ^ x248;
  assign n7360 = ~n5442 & n7359;
  assign n7361 = n7360 ^ x248;
  assign n7362 = x577 ^ x238;
  assign n7363 = ~n5429 & n7362;
  assign n7364 = n7363 ^ x238;
  assign n7365 = x578 ^ x249;
  assign n7366 = ~n5282 & n7365;
  assign n7367 = n7366 ^ x249;
  assign n7368 = x579 ^ x249;
  assign n7369 = ~n5274 & n7368;
  assign n7370 = n7369 ^ x249;
  assign n7371 = x580 ^ x245;
  assign n7372 = ~n5429 & n7371;
  assign n7373 = n7372 ^ x245;
  assign n7374 = x581 ^ x235;
  assign n7375 = ~n5282 & n7374;
  assign n7376 = n7375 ^ x235;
  assign n7377 = x582 ^ x240;
  assign n7378 = ~n5282 & n7377;
  assign n7379 = n7378 ^ x240;
  assign n7380 = x584 ^ x245;
  assign n7381 = ~n5282 & n7380;
  assign n7382 = n7381 ^ x245;
  assign n7383 = x585 ^ x244;
  assign n7384 = ~n5282 & n7383;
  assign n7385 = n7384 ^ x244;
  assign n7386 = x586 ^ x242;
  assign n7387 = ~n5282 & n7386;
  assign n7388 = n7387 ^ x242;
  assign n7389 = n4580 ^ x587;
  assign n7390 = x230 & n7389;
  assign n7391 = n7390 ^ x587;
  assign n7392 = ~x123 & x824;
  assign n7393 = x950 & n7392;
  assign n7394 = n7393 ^ x591;
  assign n7395 = n7394 ^ x591;
  assign n7396 = x591 ^ x588;
  assign n7397 = ~n7395 & n7396;
  assign n7398 = n7397 ^ x591;
  assign n7399 = n6574 & n7398;
  assign n7403 = x237 ^ x206;
  assign n7404 = n7403 ^ x206;
  assign n7405 = x206 ^ x204;
  assign n7406 = n7404 & n7405;
  assign n7407 = n7406 ^ x206;
  assign n7400 = x218 ^ x205;
  assign n7401 = ~x237 & n7400;
  assign n7402 = n7401 ^ x205;
  assign n7408 = n7407 ^ n7402;
  assign n7409 = x233 & n7408;
  assign n7410 = n7409 ^ n7402;
  assign n7411 = n5298 & ~n7410;
  assign n7415 = x237 ^ x220;
  assign n7416 = n7415 ^ x220;
  assign n7417 = x220 ^ x201;
  assign n7418 = n7416 & n7417;
  assign n7419 = n7418 ^ x220;
  assign n7412 = x203 ^ x202;
  assign n7413 = ~x237 & n7412;
  assign n7414 = n7413 ^ x202;
  assign n7420 = n7419 ^ n7414;
  assign n7421 = x233 & n7420;
  assign n7422 = n7421 ^ n7414;
  assign n7423 = n5267 & ~n7422;
  assign n7424 = ~n7411 & ~n7423;
  assign n7425 = x590 ^ x588;
  assign n7426 = n7393 ^ x590;
  assign n7427 = n7426 ^ x590;
  assign n7428 = n7425 & n7427;
  assign n7429 = n7428 ^ x590;
  assign n7430 = n6574 & ~n7429;
  assign n7431 = x592 ^ x591;
  assign n7432 = n7393 ^ x592;
  assign n7433 = n7432 ^ x592;
  assign n7434 = n7431 & ~n7433;
  assign n7435 = n7434 ^ x592;
  assign n7436 = n6574 & n7435;
  assign n7437 = x592 ^ x590;
  assign n7438 = n7433 & n7437;
  assign n7439 = n7438 ^ x592;
  assign n7440 = n6574 & n7439;
  assign n7480 = x248 & ~x554;
  assign n7481 = ~x247 & x552;
  assign n7482 = ~n7480 & ~n7481;
  assign n7483 = ~x240 & x551;
  assign n7484 = ~n7088 & ~n7483;
  assign n7485 = n7482 & n7484;
  assign n7486 = ~x233 & ~n7079;
  assign n7487 = n7485 & n7486;
  assign n7488 = x240 & ~x551;
  assign n7489 = ~x248 & x554;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = x247 & ~x552;
  assign n7492 = n7490 & ~n7491;
  assign n7493 = n7487 & n7492;
  assign n7494 = ~n7310 & ~n7362;
  assign n7495 = ~n7076 & ~n7371;
  assign n7496 = n7494 & n7495;
  assign n7497 = ~n7268 & ~n7286;
  assign n7498 = n7271 & ~n7280;
  assign n7499 = n7497 & n7498;
  assign n7500 = n7496 & n7499;
  assign n7501 = n7493 & n7500;
  assign n7502 = ~x241 & x490;
  assign n7503 = x233 & ~n7502;
  assign n7504 = ~n7262 & n7503;
  assign n7505 = ~n7070 & ~n7256;
  assign n7506 = n7504 & n7505;
  assign n7507 = x241 & ~x490;
  assign n7508 = ~n7094 & ~n7507;
  assign n7509 = n7506 & n7508;
  assign n7510 = ~n7073 & ~n7259;
  assign n7511 = ~n7100 & ~n7265;
  assign n7512 = n7510 & n7511;
  assign n7513 = ~n7097 & ~n7253;
  assign n7514 = n7103 & ~n7106;
  assign n7515 = n7513 & n7514;
  assign n7516 = n7512 & n7515;
  assign n7517 = n7509 & n7516;
  assign n7518 = ~n7501 & ~n7517;
  assign n7441 = ~x238 & x507;
  assign n7442 = x233 & ~n7441;
  assign n7443 = ~n7235 & n7442;
  assign n7444 = ~n7133 & ~n7220;
  assign n7445 = n7443 & n7444;
  assign n7446 = x238 & ~x507;
  assign n7447 = ~n7145 & ~n7446;
  assign n7448 = n7445 & n7447;
  assign n7449 = ~n7226 & ~n7292;
  assign n7450 = ~n7139 & ~n7295;
  assign n7451 = n7449 & n7450;
  assign n7452 = ~n7148 & ~n7232;
  assign n7453 = n7223 & ~n7229;
  assign n7454 = n7452 & n7453;
  assign n7455 = n7451 & n7454;
  assign n7456 = n7448 & n7455;
  assign n7457 = ~x245 & x503;
  assign n7458 = ~x246 & x499;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = x241 & ~x500;
  assign n7461 = ~n7238 & ~n7460;
  assign n7462 = n7459 & n7461;
  assign n7463 = ~x233 & ~n7109;
  assign n7464 = n7462 & n7463;
  assign n7465 = x246 & ~x499;
  assign n7466 = ~x241 & x500;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = x245 & ~x503;
  assign n7469 = n7467 & ~n7468;
  assign n7470 = n7464 & n7469;
  assign n7471 = ~n7124 & ~n7250;
  assign n7472 = ~n7127 & ~n7241;
  assign n7473 = n7471 & n7472;
  assign n7474 = ~n7136 & ~n7244;
  assign n7475 = n7112 & ~n7247;
  assign n7476 = n7474 & n7475;
  assign n7477 = n7473 & n7476;
  assign n7478 = n7470 & n7477;
  assign n7479 = ~n7456 & ~n7478;
  assign n7519 = n7518 ^ n7479;
  assign n7520 = ~x237 & n7519;
  assign n7521 = n7520 ^ n7479;
  assign n7522 = n5298 & ~n7521;
  assign n7523 = ~x245 & x514;
  assign n7524 = ~n7368 & ~n7523;
  assign n7525 = x233 & n7524;
  assign n7526 = ~n7169 & ~n7298;
  assign n7527 = n7525 & n7526;
  assign n7528 = x245 & ~x514;
  assign n7529 = ~n7064 & ~n7528;
  assign n7530 = n7527 & n7529;
  assign n7531 = ~n7154 & ~n7160;
  assign n7532 = ~n7151 & ~n7166;
  assign n7533 = n7531 & n7532;
  assign n7534 = n7085 & ~n7157;
  assign n7535 = ~n7082 & ~n7172;
  assign n7536 = n7534 & n7535;
  assign n7537 = n7533 & n7536;
  assign n7538 = n7530 & n7537;
  assign n7539 = x237 & ~n7538;
  assign n7540 = ~x248 & x521;
  assign n7541 = ~x233 & ~n7540;
  assign n7542 = ~n7353 & n7541;
  assign n7543 = ~n7187 & ~n7365;
  assign n7544 = n7542 & n7543;
  assign n7545 = x248 & ~x521;
  assign n7546 = ~n7383 & ~n7545;
  assign n7547 = n7544 & n7546;
  assign n7548 = n7178 & ~n7380;
  assign n7549 = ~n7175 & ~n7181;
  assign n7550 = n7548 & n7549;
  assign n7551 = ~n7304 & ~n7386;
  assign n7552 = ~n7374 & ~n7377;
  assign n7553 = n7551 & n7552;
  assign n7554 = n7550 & n7553;
  assign n7555 = n7547 & n7554;
  assign n7556 = n7539 & ~n7555;
  assign n7557 = n5267 & ~n7556;
  assign n7558 = n7193 & ~n7196;
  assign n7559 = ~n7205 & ~n7208;
  assign n7560 = n7558 & n7559;
  assign n7561 = ~n7199 & ~n7356;
  assign n7562 = ~n7190 & ~n7350;
  assign n7563 = n7561 & n7562;
  assign n7564 = n7560 & n7563;
  assign n7565 = ~x244 & x572;
  assign n7566 = ~x247 & x527;
  assign n7567 = ~n7565 & ~n7566;
  assign n7568 = ~n7359 & n7567;
  assign n7569 = x247 & ~x527;
  assign n7570 = x233 & ~n7569;
  assign n7571 = ~n7344 & n7570;
  assign n7572 = n7568 & n7571;
  assign n7573 = n7564 & n7572;
  assign n7574 = x244 & ~x572;
  assign n7575 = ~n7211 & ~n7574;
  assign n7576 = n7573 & n7575;
  assign n7577 = ~n7316 & ~n7341;
  assign n7578 = ~n7301 & ~n7313;
  assign n7579 = n7577 & n7578;
  assign n7580 = ~n7217 & ~n7335;
  assign n7581 = ~n7115 & n7338;
  assign n7582 = n7580 & n7581;
  assign n7583 = n7579 & n7582;
  assign n7584 = ~x249 & x482;
  assign n7585 = ~x233 & ~n7584;
  assign n7586 = ~n7307 & n7585;
  assign n7587 = ~n7214 & ~n7319;
  assign n7588 = n7586 & n7587;
  assign n7589 = n7583 & n7588;
  assign n7590 = x249 & ~x482;
  assign n7591 = ~n7289 & ~n7590;
  assign n7592 = n7589 & n7591;
  assign n7593 = ~n7576 & ~n7592;
  assign n7594 = ~x237 & n7593;
  assign n7595 = n7557 & ~n7594;
  assign n7596 = ~n7522 & ~n7595;
  assign n7597 = ~x806 & x990;
  assign n7598 = x600 & n7597;
  assign n7599 = n7598 ^ x594;
  assign n7600 = ~x332 & n7599;
  assign n7601 = x605 & ~x806;
  assign n7602 = n6970 & n7601;
  assign n7603 = n7602 ^ x595;
  assign n7604 = ~x332 & n7603;
  assign n7605 = n6968 & n7597;
  assign n7606 = x595 & x597;
  assign n7607 = n7605 & n7606;
  assign n7608 = n7607 ^ x596;
  assign n7609 = ~x332 & n7608;
  assign n7610 = n7605 ^ x597;
  assign n7611 = ~x332 & n7610;
  assign n7612 = ~x882 & n1571;
  assign n7613 = x947 & n7612;
  assign n7614 = x598 & ~n7613;
  assign n7615 = x740 & x780;
  assign n7616 = n2349 & n7615;
  assign n7617 = ~n7614 & ~n7616;
  assign n7618 = x596 & n7607;
  assign n7619 = n7618 ^ x599;
  assign n7620 = ~x332 & n7619;
  assign n7621 = n7597 ^ x600;
  assign n7622 = ~x332 & n7621;
  assign n7623 = x806 ^ x601;
  assign n7624 = n7623 ^ x601;
  assign n7625 = x989 ^ x601;
  assign n7626 = ~n7624 & n7625;
  assign n7627 = n7626 ^ x601;
  assign n7628 = ~x332 & n7627;
  assign n7629 = n4606 ^ x602;
  assign n7630 = x230 & n7629;
  assign n7631 = n7630 ^ x602;
  assign n7632 = x832 & ~x980;
  assign n7633 = x1060 & n7632;
  assign n7634 = x1038 & ~x1061;
  assign n7635 = n7633 & n7634;
  assign n7636 = x952 & n7635;
  assign n7637 = n7636 ^ x603;
  assign n7638 = n7637 ^ x603;
  assign n7639 = x1100 ^ x603;
  assign n7640 = n7638 & n7639;
  assign n7641 = n7640 ^ x603;
  assign n7642 = n7641 ^ x872;
  assign n7643 = n7642 ^ n7641;
  assign n7644 = n7641 ^ x871;
  assign n7645 = n7644 ^ n7641;
  assign n7646 = ~n7643 & ~n7645;
  assign n7647 = n7646 ^ n7641;
  assign n7648 = x966 & ~n7647;
  assign n7649 = n7648 ^ n7641;
  assign n7650 = x823 & n2351;
  assign n7651 = ~x299 & x983;
  assign n7652 = x907 & n7651;
  assign n7653 = x604 & ~n7652;
  assign n7654 = n7653 ^ x779;
  assign n7655 = ~n7650 & ~n7654;
  assign n7656 = n7655 ^ x779;
  assign n7657 = x806 ^ x605;
  assign n7658 = ~x332 & ~n7657;
  assign n7659 = x837 ^ x606;
  assign n7660 = n7659 ^ x1104;
  assign n7661 = n7660 ^ x606;
  assign n7662 = n7661 ^ n7659;
  assign n7663 = n7659 ^ n7636;
  assign n7664 = n7663 ^ n7659;
  assign n7665 = n7662 & n7664;
  assign n7666 = n7665 ^ n7659;
  assign n7667 = ~x966 & n7666;
  assign n7668 = n7667 ^ x837;
  assign n7669 = n7636 ^ x607;
  assign n7670 = n7669 ^ x607;
  assign n7671 = x1107 ^ x607;
  assign n7672 = n7670 & n7671;
  assign n7673 = n7672 ^ x607;
  assign n7674 = ~x966 & n7673;
  assign n7675 = n7636 ^ x608;
  assign n7676 = n7675 ^ x608;
  assign n7677 = x1116 ^ x608;
  assign n7678 = n7676 & n7677;
  assign n7679 = n7678 ^ x608;
  assign n7680 = ~x966 & n7679;
  assign n7681 = n7636 ^ x609;
  assign n7682 = n7681 ^ x609;
  assign n7683 = x1118 ^ x609;
  assign n7684 = n7682 & n7683;
  assign n7685 = n7684 ^ x609;
  assign n7686 = ~x966 & n7685;
  assign n7687 = n7636 ^ x610;
  assign n7688 = n7687 ^ x610;
  assign n7689 = x1113 ^ x610;
  assign n7690 = n7688 & n7689;
  assign n7691 = n7690 ^ x610;
  assign n7692 = ~x966 & n7691;
  assign n7693 = n7636 ^ x611;
  assign n7694 = n7693 ^ x611;
  assign n7695 = x1114 ^ x611;
  assign n7696 = n7694 & n7695;
  assign n7697 = n7696 ^ x611;
  assign n7698 = ~x966 & n7697;
  assign n7699 = n7636 ^ x612;
  assign n7700 = n7699 ^ x612;
  assign n7701 = x1111 ^ x612;
  assign n7702 = n7700 & n7701;
  assign n7703 = n7702 ^ x612;
  assign n7704 = ~x966 & n7703;
  assign n7705 = n7636 ^ x613;
  assign n7706 = n7705 ^ x613;
  assign n7707 = x1115 ^ x613;
  assign n7708 = n7706 & n7707;
  assign n7709 = n7708 ^ x613;
  assign n7710 = ~x966 & n7709;
  assign n7711 = x1102 ^ x614;
  assign n7712 = n7636 & n7711;
  assign n7713 = n7712 ^ x614;
  assign n7714 = n7713 ^ x871;
  assign n7715 = ~x966 & n7714;
  assign n7716 = n7715 ^ x871;
  assign n7717 = x907 & n7612;
  assign n7718 = ~x615 & ~n7717;
  assign n7719 = x779 & x797;
  assign n7720 = n2352 & n7719;
  assign n7721 = ~n7718 & ~n7720;
  assign n7722 = x872 ^ x616;
  assign n7723 = n7722 ^ x1101;
  assign n7724 = n7723 ^ x616;
  assign n7725 = n7724 ^ n7722;
  assign n7726 = n7722 ^ n7636;
  assign n7727 = n7726 ^ n7722;
  assign n7728 = n7725 & n7727;
  assign n7729 = n7728 ^ n7722;
  assign n7730 = ~x966 & n7729;
  assign n7731 = n7730 ^ x872;
  assign n7732 = x850 ^ x617;
  assign n7733 = n7732 ^ x1105;
  assign n7734 = n7733 ^ x617;
  assign n7735 = n7734 ^ n7732;
  assign n7736 = n7732 ^ n7636;
  assign n7737 = n7736 ^ n7732;
  assign n7738 = n7735 & n7737;
  assign n7739 = n7738 ^ n7732;
  assign n7740 = ~x966 & n7739;
  assign n7741 = n7740 ^ x850;
  assign n7742 = n7636 ^ x618;
  assign n7743 = n7742 ^ x618;
  assign n7744 = x1117 ^ x618;
  assign n7745 = n7743 & n7744;
  assign n7746 = n7745 ^ x618;
  assign n7747 = ~x966 & n7746;
  assign n7748 = n7636 ^ x619;
  assign n7749 = n7748 ^ x619;
  assign n7750 = x1122 ^ x619;
  assign n7751 = n7749 & n7750;
  assign n7752 = n7751 ^ x619;
  assign n7753 = ~x966 & n7752;
  assign n7754 = n7636 ^ x620;
  assign n7755 = n7754 ^ x620;
  assign n7756 = x1112 ^ x620;
  assign n7757 = n7755 & n7756;
  assign n7758 = n7757 ^ x620;
  assign n7759 = ~x966 & n7758;
  assign n7760 = n7636 ^ x621;
  assign n7761 = n7760 ^ x621;
  assign n7762 = x1108 ^ x621;
  assign n7763 = n7761 & n7762;
  assign n7764 = n7763 ^ x621;
  assign n7765 = ~x966 & n7764;
  assign n7766 = n7636 ^ x622;
  assign n7767 = n7766 ^ x622;
  assign n7768 = x1109 ^ x622;
  assign n7769 = n7767 & n7768;
  assign n7770 = n7769 ^ x622;
  assign n7771 = ~x966 & n7770;
  assign n7772 = n7636 ^ x623;
  assign n7773 = n7772 ^ x623;
  assign n7774 = x1106 ^ x623;
  assign n7775 = n7773 & n7774;
  assign n7776 = n7775 ^ x623;
  assign n7777 = ~x966 & n7776;
  assign n7778 = x831 & n2348;
  assign n7779 = x947 & n7651;
  assign n7780 = x624 & ~n7779;
  assign n7781 = n7780 ^ x780;
  assign n7782 = ~n7778 & ~n7781;
  assign n7783 = n7782 ^ x780;
  assign n7784 = x1066 & x1088;
  assign n7785 = ~x973 & ~x1054;
  assign n7786 = n7784 & n7785;
  assign n7787 = x832 & n7786;
  assign n7788 = ~x953 & n7787;
  assign n7789 = n7788 ^ x625;
  assign n7790 = n7789 ^ x625;
  assign n7791 = x1116 ^ x625;
  assign n7792 = n7790 & n7791;
  assign n7793 = n7792 ^ x625;
  assign n7794 = ~x962 & n7793;
  assign n7795 = n7636 ^ x626;
  assign n7796 = n7795 ^ x626;
  assign n7797 = x1121 ^ x626;
  assign n7798 = n7796 & n7797;
  assign n7799 = n7798 ^ x626;
  assign n7800 = ~x966 & n7799;
  assign n7801 = n7788 ^ x627;
  assign n7802 = n7801 ^ x627;
  assign n7803 = x1117 ^ x627;
  assign n7804 = n7802 & n7803;
  assign n7805 = n7804 ^ x627;
  assign n7806 = ~x962 & n7805;
  assign n7807 = n7788 ^ x628;
  assign n7808 = n7807 ^ x628;
  assign n7809 = x1119 ^ x628;
  assign n7810 = n7808 & n7809;
  assign n7811 = n7810 ^ x628;
  assign n7812 = ~x962 & n7811;
  assign n7813 = n7636 ^ x629;
  assign n7814 = n7813 ^ x629;
  assign n7815 = x1119 ^ x629;
  assign n7816 = n7814 & n7815;
  assign n7817 = n7816 ^ x629;
  assign n7818 = ~x966 & n7817;
  assign n7819 = n7636 ^ x630;
  assign n7820 = n7819 ^ x630;
  assign n7821 = x1120 ^ x630;
  assign n7822 = n7820 & n7821;
  assign n7823 = n7822 ^ x630;
  assign n7824 = ~x966 & n7823;
  assign n7825 = n7788 ^ x631;
  assign n7826 = n7825 ^ x631;
  assign n7827 = x1113 ^ x631;
  assign n7828 = n7826 & ~n7827;
  assign n7829 = n7828 ^ x631;
  assign n7830 = ~x962 & ~n7829;
  assign n7831 = n7788 ^ x632;
  assign n7832 = n7831 ^ x632;
  assign n7833 = x1115 ^ x632;
  assign n7834 = n7832 & ~n7833;
  assign n7835 = n7834 ^ x632;
  assign n7836 = ~x962 & ~n7835;
  assign n7837 = n7636 ^ x633;
  assign n7838 = n7837 ^ x633;
  assign n7839 = x1110 ^ x633;
  assign n7840 = n7838 & n7839;
  assign n7841 = n7840 ^ x633;
  assign n7842 = ~x966 & n7841;
  assign n7843 = n7788 ^ x634;
  assign n7844 = n7843 ^ x634;
  assign n7845 = x1110 ^ x634;
  assign n7846 = n7844 & n7845;
  assign n7847 = n7846 ^ x634;
  assign n7848 = ~x962 & n7847;
  assign n7849 = n7788 ^ x635;
  assign n7850 = n7849 ^ x635;
  assign n7851 = x1112 ^ x635;
  assign n7852 = n7850 & ~n7851;
  assign n7853 = n7852 ^ x635;
  assign n7854 = ~x962 & ~n7853;
  assign n7855 = n7636 ^ x636;
  assign n7856 = n7855 ^ x636;
  assign n7857 = x1127 ^ x636;
  assign n7858 = n7856 & n7857;
  assign n7859 = n7858 ^ x636;
  assign n7860 = ~x966 & n7859;
  assign n7861 = n7788 ^ x637;
  assign n7862 = n7861 ^ x637;
  assign n7863 = x1105 ^ x637;
  assign n7864 = n7862 & n7863;
  assign n7865 = n7864 ^ x637;
  assign n7866 = ~x962 & n7865;
  assign n7867 = n7788 ^ x638;
  assign n7868 = n7867 ^ x638;
  assign n7869 = x1107 ^ x638;
  assign n7870 = n7868 & n7869;
  assign n7871 = n7870 ^ x638;
  assign n7872 = ~x962 & n7871;
  assign n7873 = n7788 ^ x639;
  assign n7874 = n7873 ^ x639;
  assign n7875 = x1109 ^ x639;
  assign n7876 = n7874 & n7875;
  assign n7877 = n7876 ^ x639;
  assign n7878 = ~x962 & n7877;
  assign n7879 = n7636 ^ x640;
  assign n7880 = n7879 ^ x640;
  assign n7881 = x1128 ^ x640;
  assign n7882 = n7880 & n7881;
  assign n7883 = n7882 ^ x640;
  assign n7884 = ~x966 & n7883;
  assign n7885 = n7788 ^ x641;
  assign n7886 = n7885 ^ x641;
  assign n7887 = x1121 ^ x641;
  assign n7888 = n7886 & n7887;
  assign n7889 = n7888 ^ x641;
  assign n7890 = ~x962 & n7889;
  assign n7891 = n7636 ^ x642;
  assign n7892 = n7891 ^ x642;
  assign n7893 = x1103 ^ x642;
  assign n7894 = n7892 & n7893;
  assign n7895 = n7894 ^ x642;
  assign n7896 = ~x966 & n7895;
  assign n7897 = n7788 ^ x643;
  assign n7898 = n7897 ^ x643;
  assign n7899 = x1104 ^ x643;
  assign n7900 = n7898 & n7899;
  assign n7901 = n7900 ^ x643;
  assign n7902 = ~x962 & n7901;
  assign n7903 = n7636 ^ x644;
  assign n7904 = n7903 ^ x644;
  assign n7905 = x1123 ^ x644;
  assign n7906 = n7904 & n7905;
  assign n7907 = n7906 ^ x644;
  assign n7908 = ~x966 & n7907;
  assign n7909 = n7636 ^ x645;
  assign n7910 = n7909 ^ x645;
  assign n7911 = x1125 ^ x645;
  assign n7912 = n7910 & n7911;
  assign n7913 = n7912 ^ x645;
  assign n7914 = ~x966 & n7913;
  assign n7915 = n7788 ^ x646;
  assign n7916 = n7915 ^ x646;
  assign n7917 = x1114 ^ x646;
  assign n7918 = n7916 & ~n7917;
  assign n7919 = n7918 ^ x646;
  assign n7920 = ~x962 & ~n7919;
  assign n7921 = n7788 ^ x647;
  assign n7922 = n7921 ^ x647;
  assign n7923 = x1120 ^ x647;
  assign n7924 = n7922 & n7923;
  assign n7925 = n7924 ^ x647;
  assign n7926 = ~x962 & n7925;
  assign n7927 = n7788 ^ x648;
  assign n7928 = n7927 ^ x648;
  assign n7929 = x1122 ^ x648;
  assign n7930 = n7928 & n7929;
  assign n7931 = n7930 ^ x648;
  assign n7932 = ~x962 & n7931;
  assign n7933 = n7788 ^ x649;
  assign n7934 = n7933 ^ x649;
  assign n7935 = x1126 ^ x649;
  assign n7936 = n7934 & ~n7935;
  assign n7937 = n7936 ^ x649;
  assign n7938 = ~x962 & ~n7937;
  assign n7939 = n7788 ^ x650;
  assign n7940 = n7939 ^ x650;
  assign n7941 = x1127 ^ x650;
  assign n7942 = n7940 & ~n7941;
  assign n7943 = n7942 ^ x650;
  assign n7944 = ~x962 & ~n7943;
  assign n7945 = n7636 ^ x651;
  assign n7946 = n7945 ^ x651;
  assign n7947 = x1130 ^ x651;
  assign n7948 = n7946 & n7947;
  assign n7949 = n7948 ^ x651;
  assign n7950 = ~x966 & n7949;
  assign n7951 = n7636 ^ x652;
  assign n7952 = n7951 ^ x652;
  assign n7953 = x1131 ^ x652;
  assign n7954 = n7952 & n7953;
  assign n7955 = n7954 ^ x652;
  assign n7956 = ~x966 & n7955;
  assign n7957 = n7636 ^ x653;
  assign n7958 = n7957 ^ x653;
  assign n7959 = x1129 ^ x653;
  assign n7960 = n7958 & n7959;
  assign n7961 = n7960 ^ x653;
  assign n7962 = ~x966 & n7961;
  assign n7963 = n7788 ^ x654;
  assign n7964 = n7963 ^ x654;
  assign n7965 = x1130 ^ x654;
  assign n7966 = n7964 & ~n7965;
  assign n7967 = n7966 ^ x654;
  assign n7968 = ~x962 & ~n7967;
  assign n7969 = n7788 ^ x655;
  assign n7970 = n7969 ^ x655;
  assign n7971 = x1124 ^ x655;
  assign n7972 = n7970 & ~n7971;
  assign n7973 = n7972 ^ x655;
  assign n7974 = ~x962 & ~n7973;
  assign n7975 = n7636 ^ x656;
  assign n7976 = n7975 ^ x656;
  assign n7977 = x1126 ^ x656;
  assign n7978 = n7976 & n7977;
  assign n7979 = n7978 ^ x656;
  assign n7980 = ~x966 & n7979;
  assign n7981 = n7788 ^ x657;
  assign n7982 = n7981 ^ x657;
  assign n7983 = x1131 ^ x657;
  assign n7984 = n7982 & ~n7983;
  assign n7985 = n7984 ^ x657;
  assign n7986 = ~x962 & ~n7985;
  assign n7987 = n7636 ^ x658;
  assign n7988 = n7987 ^ x658;
  assign n7989 = x1124 ^ x658;
  assign n7990 = n7988 & n7989;
  assign n7991 = n7990 ^ x658;
  assign n7992 = ~x966 & n7991;
  assign n7993 = x266 & x992;
  assign n7994 = ~x280 & n7993;
  assign n7995 = ~x269 & n7994;
  assign n7996 = ~x281 & ~x282;
  assign n7997 = n7995 & n7996;
  assign n7998 = ~x270 & ~x277;
  assign n7999 = ~x264 & n7998;
  assign n8000 = n7997 & n7999;
  assign n8001 = ~x265 & n8000;
  assign n8002 = n8001 ^ x274;
  assign n8003 = n7788 ^ x660;
  assign n8004 = n8003 ^ x660;
  assign n8005 = x1118 ^ x660;
  assign n8006 = n8004 & n8005;
  assign n8007 = n8006 ^ x660;
  assign n8008 = ~x962 & n8007;
  assign n8009 = n7788 ^ x661;
  assign n8010 = n8009 ^ x661;
  assign n8011 = x1101 ^ x661;
  assign n8012 = n8010 & n8011;
  assign n8013 = n8012 ^ x661;
  assign n8014 = ~x962 & n8013;
  assign n8015 = n7788 ^ x662;
  assign n8016 = n8015 ^ x662;
  assign n8017 = x1102 ^ x662;
  assign n8018 = n8016 & n8017;
  assign n8019 = n8018 ^ x662;
  assign n8020 = ~x962 & n8019;
  assign n8021 = x592 ^ x365;
  assign n8022 = n8021 ^ x365;
  assign n8023 = x365 ^ x334;
  assign n8024 = ~n8022 & n8023;
  assign n8025 = n8024 ^ x365;
  assign n8026 = n7431 & n8025;
  assign n8027 = n3754 & n8026;
  assign n8028 = x588 & n2809;
  assign n8029 = x464 & n8028;
  assign n8030 = ~n8027 & ~n8029;
  assign n8031 = n1536 & n8030;
  assign n8032 = ~x588 & ~n2809;
  assign n8033 = n2806 & n8032;
  assign n8034 = x323 & n8033;
  assign n8035 = n8031 & ~n8034;
  assign n8036 = x1065 ^ x257;
  assign n8037 = x199 & n8036;
  assign n8038 = n8037 ^ x257;
  assign n8039 = ~n1536 & ~n8038;
  assign n8040 = n2872 & ~n8039;
  assign n8041 = ~n8035 & n8040;
  assign n8042 = ~x1137 & ~x1138;
  assign n8043 = ~n2872 & n8042;
  assign n8047 = x855 ^ x766;
  assign n8048 = ~x1136 & n8047;
  assign n8049 = n8048 ^ x766;
  assign n8044 = x815 ^ x633;
  assign n8045 = ~x1136 & n8044;
  assign n8046 = n8045 ^ x633;
  assign n8050 = n8049 ^ n8046;
  assign n8051 = x1134 & n8050;
  assign n8052 = n8051 ^ n8046;
  assign n8053 = n8052 ^ x1135;
  assign n8054 = n8053 ^ n8052;
  assign n8055 = x784 ^ x634;
  assign n8056 = ~x1136 & n8055;
  assign n8057 = n8056 ^ x634;
  assign n8058 = n8057 ^ x1134;
  assign n8059 = n8058 ^ n8057;
  assign n8060 = n8059 ^ x1135;
  assign n8061 = x1136 ^ x700;
  assign n8062 = x1136 & n8061;
  assign n8063 = n8062 ^ n8057;
  assign n8064 = n8063 ^ x1136;
  assign n8065 = n8060 & n8064;
  assign n8066 = n8065 ^ n8062;
  assign n8067 = n8066 ^ x1136;
  assign n8068 = n8067 ^ n8052;
  assign n8069 = n8054 & n8068;
  assign n8070 = n8069 ^ n8052;
  assign n8071 = n8043 & n8070;
  assign n8072 = ~n8041 & ~n8071;
  assign n8073 = x592 ^ x404;
  assign n8074 = n8073 ^ x404;
  assign n8075 = x404 ^ x380;
  assign n8076 = n8074 & n8075;
  assign n8077 = n8076 ^ x404;
  assign n8078 = n7431 & n8077;
  assign n8079 = n3754 & n8078;
  assign n8080 = x429 & n8028;
  assign n8081 = ~n8079 & ~n8080;
  assign n8082 = n1536 & n8081;
  assign n8083 = x355 & n8033;
  assign n8084 = n8082 & ~n8083;
  assign n8085 = x199 & n6429;
  assign n8086 = n8085 ^ x292;
  assign n8087 = ~n1536 & ~n8086;
  assign n8088 = n2872 & ~n8087;
  assign n8089 = ~n8084 & n8088;
  assign n8093 = x872 ^ x772;
  assign n8094 = ~x1136 & n8093;
  assign n8095 = n8094 ^ x772;
  assign n8090 = x811 ^ x614;
  assign n8091 = ~x1136 & n8090;
  assign n8092 = n8091 ^ x614;
  assign n8096 = n8095 ^ n8092;
  assign n8097 = x1134 & n8096;
  assign n8098 = n8097 ^ n8092;
  assign n8099 = n8098 ^ x1135;
  assign n8100 = n8099 ^ n8098;
  assign n8101 = x785 ^ x662;
  assign n8102 = ~x1136 & n8101;
  assign n8103 = n8102 ^ x662;
  assign n8104 = n8103 ^ x1134;
  assign n8105 = n8104 ^ n8103;
  assign n8106 = n8105 ^ x1135;
  assign n8107 = x1136 ^ x727;
  assign n8108 = x1136 & n8107;
  assign n8109 = n8108 ^ n8103;
  assign n8110 = n8109 ^ x1136;
  assign n8111 = n8106 & n8110;
  assign n8112 = n8111 ^ n8108;
  assign n8113 = n8112 ^ x1136;
  assign n8114 = n8113 ^ n8098;
  assign n8115 = n8100 & n8114;
  assign n8116 = n8115 ^ n8098;
  assign n8117 = n8043 & n8116;
  assign n8118 = ~n8089 & ~n8117;
  assign n8119 = n7788 ^ x665;
  assign n8120 = n8119 ^ x665;
  assign n8121 = x1108 ^ x665;
  assign n8122 = n8120 & n8121;
  assign n8123 = n8122 ^ x665;
  assign n8124 = ~x962 & n8123;
  assign n8125 = x592 ^ x456;
  assign n8126 = n8125 ^ x456;
  assign n8127 = x456 ^ x337;
  assign n8128 = n8126 & n8127;
  assign n8129 = n8128 ^ x456;
  assign n8130 = n7431 & n8129;
  assign n8131 = n3754 & n8130;
  assign n8132 = x443 & n8028;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = n1536 & n8133;
  assign n8135 = x441 & n8033;
  assign n8136 = n8134 & ~n8135;
  assign n8137 = x199 & n6444;
  assign n8138 = n8137 ^ x297;
  assign n8139 = ~n1536 & ~n8138;
  assign n8140 = n2872 & ~n8139;
  assign n8141 = ~n8136 & n8140;
  assign n8145 = x1136 ^ x873;
  assign n8146 = n8145 ^ x873;
  assign n8147 = x873 ^ x764;
  assign n8148 = n8146 & n8147;
  assign n8149 = n8148 ^ x873;
  assign n8142 = x799 ^ x607;
  assign n8143 = ~x1136 & ~n8142;
  assign n8144 = n8143 ^ x607;
  assign n8150 = n8149 ^ n8144;
  assign n8151 = x1134 & n8150;
  assign n8152 = n8151 ^ n8144;
  assign n8153 = n8152 ^ x1135;
  assign n8154 = n8153 ^ n8152;
  assign n8155 = x790 ^ x638;
  assign n8156 = ~x1136 & n8155;
  assign n8157 = n8156 ^ x638;
  assign n8158 = n8157 ^ x1134;
  assign n8159 = n8158 ^ n8157;
  assign n8160 = n8159 ^ x1135;
  assign n8161 = x1136 ^ x691;
  assign n8162 = x1136 & n8161;
  assign n8163 = n8162 ^ n8157;
  assign n8164 = n8163 ^ x1136;
  assign n8165 = n8160 & n8164;
  assign n8166 = n8165 ^ n8162;
  assign n8167 = n8166 ^ x1136;
  assign n8168 = n8167 ^ n8152;
  assign n8169 = n8154 & n8168;
  assign n8170 = n8169 ^ n8152;
  assign n8171 = n8043 & n8170;
  assign n8172 = ~n8141 & ~n8171;
  assign n8202 = x458 & n8033;
  assign n8203 = x592 ^ x338;
  assign n8204 = n8203 ^ x338;
  assign n8205 = x338 ^ x319;
  assign n8206 = ~n8204 & n8205;
  assign n8207 = n8206 ^ x338;
  assign n8208 = n7431 & n8207;
  assign n8209 = n3754 & n8208;
  assign n8210 = x444 & n8028;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = ~n8202 & n8211;
  assign n8213 = n8212 ^ n1536;
  assign n8214 = n8213 ^ n8212;
  assign n8215 = x199 & n6435;
  assign n8216 = n8215 ^ x294;
  assign n8217 = n8216 ^ n8212;
  assign n8218 = ~n8214 & ~n8217;
  assign n8219 = n8218 ^ n8212;
  assign n8176 = x1136 ^ x871;
  assign n8177 = n8176 ^ x871;
  assign n8178 = x871 ^ x763;
  assign n8179 = n8177 & n8178;
  assign n8180 = n8179 ^ x871;
  assign n8173 = x809 ^ x642;
  assign n8174 = ~x1136 & ~n8173;
  assign n8175 = n8174 ^ x642;
  assign n8181 = n8180 ^ n8175;
  assign n8182 = x1134 & n8181;
  assign n8183 = n8182 ^ n8175;
  assign n8184 = n8183 ^ x1135;
  assign n8185 = n8184 ^ n8183;
  assign n8186 = x792 ^ x681;
  assign n8187 = ~x1136 & n8186;
  assign n8188 = n8187 ^ x681;
  assign n8189 = n8188 ^ x1134;
  assign n8190 = n8189 ^ n8188;
  assign n8191 = n8190 ^ x1135;
  assign n8192 = x1136 ^ x699;
  assign n8193 = x1136 & n8192;
  assign n8194 = n8193 ^ n8188;
  assign n8195 = n8194 ^ x1136;
  assign n8196 = n8191 & n8195;
  assign n8197 = n8196 ^ n8193;
  assign n8198 = n8197 ^ x1136;
  assign n8199 = n8198 ^ n8183;
  assign n8200 = n8185 & n8199;
  assign n8201 = n8200 ^ n8183;
  assign n8220 = n8219 ^ n8201;
  assign n8221 = n8220 ^ n8219;
  assign n8222 = n8219 ^ n8042;
  assign n8223 = n8222 ^ n8219;
  assign n8224 = n8221 & n8223;
  assign n8225 = n8224 ^ n8219;
  assign n8226 = ~n2872 & ~n8225;
  assign n8227 = n8226 ^ n8219;
  assign n8249 = x837 ^ x759;
  assign n8250 = ~x1136 & n8249;
  assign n8251 = n8250 ^ x759;
  assign n8246 = x981 ^ x603;
  assign n8247 = ~x1136 & n8246;
  assign n8248 = n8247 ^ x603;
  assign n8252 = n8251 ^ n8248;
  assign n8253 = x1134 & n8252;
  assign n8254 = n8253 ^ n8248;
  assign n8255 = n8254 ^ x1135;
  assign n8256 = n8255 ^ n8254;
  assign n8257 = x778 ^ x680;
  assign n8258 = ~x1136 & n8257;
  assign n8259 = n8258 ^ x680;
  assign n8260 = n8259 ^ x1134;
  assign n8261 = n8260 ^ n8259;
  assign n8262 = n8261 ^ x1135;
  assign n8263 = x1136 ^ x696;
  assign n8264 = x1136 & n8263;
  assign n8265 = n8264 ^ n8259;
  assign n8266 = n8265 ^ x1136;
  assign n8267 = n8262 & n8266;
  assign n8268 = n8267 ^ n8264;
  assign n8269 = n8268 ^ x1136;
  assign n8270 = n8269 ^ n8254;
  assign n8271 = n8256 & n8270;
  assign n8272 = n8271 ^ n8254;
  assign n8228 = x342 & n8033;
  assign n8229 = x592 ^ x390;
  assign n8230 = n8229 ^ x390;
  assign n8231 = x390 ^ x363;
  assign n8232 = n8230 & n8231;
  assign n8233 = n8232 ^ x390;
  assign n8234 = n7431 & n8233;
  assign n8235 = n3754 & n8234;
  assign n8236 = x414 & n8028;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = ~n8228 & n8237;
  assign n8239 = n8238 ^ n1536;
  assign n8240 = n8239 ^ n8238;
  assign n8241 = x199 & n6426;
  assign n8242 = n8241 ^ x291;
  assign n8243 = n8242 ^ n8238;
  assign n8244 = ~n8240 & ~n8243;
  assign n8245 = n8244 ^ n8238;
  assign n8273 = n8272 ^ n8245;
  assign n8274 = n8273 ^ n8245;
  assign n8275 = n8245 ^ n8042;
  assign n8276 = n8275 ^ n8245;
  assign n8277 = n8274 & n8276;
  assign n8278 = n8277 ^ n8245;
  assign n8279 = ~n2872 & ~n8278;
  assign n8280 = n8279 ^ n8245;
  assign n8281 = n7788 ^ x669;
  assign n8282 = n8281 ^ x669;
  assign n8283 = x1125 ^ x669;
  assign n8284 = n8282 & ~n8283;
  assign n8285 = n8284 ^ x669;
  assign n8286 = ~x962 & ~n8285;
  assign n8291 = x1135 ^ x695;
  assign n8292 = n8291 ^ x695;
  assign n8293 = ~n5418 & ~n8292;
  assign n8294 = n8293 ^ x695;
  assign n8287 = x1135 ^ x745;
  assign n8288 = n8287 ^ x745;
  assign n8289 = n4733 & n8288;
  assign n8290 = n8289 ^ x745;
  assign n8295 = n8294 ^ n8290;
  assign n8296 = ~x1134 & n8295;
  assign n8297 = n8296 ^ n8290;
  assign n8298 = x1136 & ~n8297;
  assign n8299 = ~x1135 & ~x1136;
  assign n8300 = x1134 & n8299;
  assign n8301 = x852 & n8300;
  assign n8302 = ~n8298 & ~n8301;
  assign n8303 = n8043 & ~n8302;
  assign n8304 = x415 & n8028;
  assign n8305 = n1536 & ~n8304;
  assign n8306 = x391 & n2703;
  assign n8307 = x364 & ~x590;
  assign n8308 = ~x591 & n8307;
  assign n8309 = ~n8306 & ~n8308;
  assign n8310 = x343 & n2806;
  assign n8311 = n8309 & ~n8310;
  assign n8312 = n8032 & ~n8311;
  assign n8313 = n8305 & ~n8312;
  assign n8314 = x1062 ^ x258;
  assign n8315 = x199 & n8314;
  assign n8316 = n8315 ^ x258;
  assign n8317 = ~n1536 & ~n8316;
  assign n8318 = n2872 & ~n8317;
  assign n8319 = ~n8313 & n8318;
  assign n8320 = ~n8303 & ~n8319;
  assign n8321 = x592 ^ x447;
  assign n8322 = n8321 ^ x447;
  assign n8323 = x447 ^ x333;
  assign n8324 = ~n8322 & n8323;
  assign n8325 = n8324 ^ x447;
  assign n8326 = n7431 & n8325;
  assign n8327 = n3754 & n8326;
  assign n8328 = x453 & n8028;
  assign n8329 = ~n8327 & ~n8328;
  assign n8330 = n1536 & n8329;
  assign n8331 = x327 & n8033;
  assign n8332 = n8330 & ~n8331;
  assign n8333 = x1040 ^ x261;
  assign n8334 = x199 & n8333;
  assign n8335 = n8334 ^ x261;
  assign n8336 = ~n1536 & ~n8335;
  assign n8337 = n2872 & ~n8336;
  assign n8338 = ~n8332 & n8337;
  assign n8343 = x1135 ^ x646;
  assign n8344 = n8343 ^ x646;
  assign n8345 = x646 ^ x611;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = n8346 ^ x646;
  assign n8339 = x1135 ^ x741;
  assign n8340 = n8339 ^ x741;
  assign n8341 = n4788 & n8340;
  assign n8342 = n8341 ^ x741;
  assign n8348 = n8347 ^ n8342;
  assign n8349 = ~x1134 & n8348;
  assign n8350 = n8349 ^ n8342;
  assign n8351 = x1136 & ~n8350;
  assign n8352 = x865 & n8300;
  assign n8353 = ~n8351 & ~n8352;
  assign n8354 = n8043 & ~n8353;
  assign n8355 = ~n8338 & ~n8354;
  assign n8383 = x320 & n8033;
  assign n8384 = x592 ^ x397;
  assign n8385 = n8384 ^ x397;
  assign n8386 = x397 ^ x372;
  assign n8387 = n8385 & n8386;
  assign n8388 = n8387 ^ x397;
  assign n8389 = n7431 & n8388;
  assign n8390 = n3754 & n8389;
  assign n8391 = x422 & n8028;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = ~n8383 & n8392;
  assign n8394 = n8393 ^ n1536;
  assign n8395 = n8394 ^ n8393;
  assign n8396 = x199 & n6423;
  assign n8397 = n8396 ^ x290;
  assign n8398 = n8397 ^ n8393;
  assign n8399 = ~n8395 & ~n8398;
  assign n8400 = n8399 ^ n8393;
  assign n8359 = x850 ^ x758;
  assign n8360 = ~x1136 & n8359;
  assign n8361 = n8360 ^ x758;
  assign n8356 = x808 ^ x616;
  assign n8357 = ~x1136 & n8356;
  assign n8358 = n8357 ^ x616;
  assign n8362 = n8361 ^ n8358;
  assign n8363 = x1134 & n8362;
  assign n8364 = n8363 ^ n8358;
  assign n8365 = n8364 ^ x1135;
  assign n8366 = n8365 ^ n8364;
  assign n8367 = x781 ^ x661;
  assign n8368 = ~x1136 & n8367;
  assign n8369 = n8368 ^ x661;
  assign n8370 = n8369 ^ x1134;
  assign n8371 = n8370 ^ n8369;
  assign n8372 = n8371 ^ x1135;
  assign n8373 = x1136 ^ x736;
  assign n8374 = x1136 & n8373;
  assign n8375 = n8374 ^ n8369;
  assign n8376 = n8375 ^ x1136;
  assign n8377 = n8372 & n8376;
  assign n8378 = n8377 ^ n8374;
  assign n8379 = n8378 ^ x1136;
  assign n8380 = n8379 ^ n8364;
  assign n8381 = n8366 & n8380;
  assign n8382 = n8381 ^ n8364;
  assign n8401 = n8400 ^ n8382;
  assign n8402 = n8401 ^ n8400;
  assign n8403 = n8400 ^ n8042;
  assign n8404 = n8403 ^ n8400;
  assign n8405 = n8402 & n8404;
  assign n8406 = n8405 ^ n8400;
  assign n8407 = ~n2872 & ~n8406;
  assign n8408 = n8407 ^ n8400;
  assign n8409 = x592 ^ x411;
  assign n8410 = n8409 ^ x411;
  assign n8411 = x411 ^ x387;
  assign n8412 = n8410 & n8411;
  assign n8413 = n8412 ^ x411;
  assign n8414 = n7431 & n8413;
  assign n8415 = n3754 & n8414;
  assign n8416 = x435 & n8028;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n1536 & n8417;
  assign n8419 = x452 & n8033;
  assign n8420 = n8418 & ~n8419;
  assign n8421 = x199 & n6438;
  assign n8422 = n8421 ^ x295;
  assign n8423 = ~n1536 & ~n8422;
  assign n8424 = n2872 & ~n8423;
  assign n8425 = ~n8420 & n8424;
  assign n8429 = x814 ^ x617;
  assign n8430 = ~x1136 & ~n8429;
  assign n8431 = n8430 ^ x617;
  assign n8426 = x866 ^ x749;
  assign n8427 = ~x1136 & n8426;
  assign n8428 = n8427 ^ x749;
  assign n8432 = n8431 ^ n8428;
  assign n8433 = ~x1134 & n8432;
  assign n8434 = n8433 ^ n8428;
  assign n8435 = n8434 ^ x1135;
  assign n8436 = n8435 ^ n8434;
  assign n8437 = x788 ^ x637;
  assign n8438 = ~x1136 & n8437;
  assign n8439 = n8438 ^ x637;
  assign n8440 = n8439 ^ x1134;
  assign n8441 = n8440 ^ n8439;
  assign n8442 = n8441 ^ x1135;
  assign n8443 = x1136 ^ x706;
  assign n8444 = x1136 & n8443;
  assign n8445 = n8444 ^ n8439;
  assign n8446 = n8445 ^ x1136;
  assign n8447 = n8442 & n8446;
  assign n8448 = n8447 ^ n8444;
  assign n8449 = n8448 ^ x1136;
  assign n8450 = n8449 ^ n8434;
  assign n8451 = n8436 & n8450;
  assign n8452 = n8451 ^ n8434;
  assign n8453 = n8043 & n8452;
  assign n8454 = ~n8425 & ~n8453;
  assign n8482 = x362 & n8033;
  assign n8483 = x592 ^ x463;
  assign n8484 = n8483 ^ x463;
  assign n8485 = x463 ^ x336;
  assign n8486 = n8484 & n8485;
  assign n8487 = n8486 ^ x463;
  assign n8488 = n7431 & n8487;
  assign n8489 = n3754 & n8488;
  assign n8490 = x437 & n8028;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = ~n8482 & n8491;
  assign n8493 = n8492 ^ n1536;
  assign n8494 = n8493 ^ n8492;
  assign n8495 = x1070 ^ x256;
  assign n8496 = x199 & n8495;
  assign n8497 = n8496 ^ x256;
  assign n8498 = n8497 ^ n8492;
  assign n8499 = ~n8494 & ~n8498;
  assign n8500 = n8499 ^ n8492;
  assign n8458 = x859 ^ x743;
  assign n8459 = ~x1136 & n8458;
  assign n8460 = n8459 ^ x743;
  assign n8455 = x804 ^ x622;
  assign n8456 = ~x1136 & n8455;
  assign n8457 = n8456 ^ x622;
  assign n8461 = n8460 ^ n8457;
  assign n8462 = x1134 & n8461;
  assign n8463 = n8462 ^ n8457;
  assign n8464 = n8463 ^ x1135;
  assign n8465 = n8464 ^ n8463;
  assign n8466 = x783 ^ x639;
  assign n8467 = ~x1136 & n8466;
  assign n8468 = n8467 ^ x639;
  assign n8469 = n8468 ^ x1134;
  assign n8470 = n8469 ^ n8468;
  assign n8471 = n8470 ^ x1135;
  assign n8472 = x1136 ^ x735;
  assign n8473 = x1136 & n8472;
  assign n8474 = n8473 ^ n8468;
  assign n8475 = n8474 ^ x1136;
  assign n8476 = n8471 & n8475;
  assign n8477 = n8476 ^ n8473;
  assign n8478 = n8477 ^ x1136;
  assign n8479 = n8478 ^ n8463;
  assign n8480 = n8465 & n8479;
  assign n8481 = n8480 ^ n8463;
  assign n8501 = n8500 ^ n8481;
  assign n8502 = n8501 ^ n8500;
  assign n8503 = n8500 ^ n8042;
  assign n8504 = n8503 ^ n8500;
  assign n8505 = n8502 & n8504;
  assign n8506 = n8505 ^ n8500;
  assign n8507 = ~n2872 & ~n8506;
  assign n8508 = n8507 ^ n8500;
  assign n8509 = x592 ^ x412;
  assign n8510 = n8509 ^ x412;
  assign n8511 = x412 ^ x388;
  assign n8512 = n8510 & n8511;
  assign n8513 = n8512 ^ x412;
  assign n8514 = n7431 & n8513;
  assign n8515 = n3754 & n8514;
  assign n8516 = x436 & n8028;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = n1536 & n8517;
  assign n8519 = x455 & n8033;
  assign n8520 = n8518 & ~n8519;
  assign n8521 = x199 & n6441;
  assign n8522 = n8521 ^ x296;
  assign n8523 = ~n1536 & ~n8522;
  assign n8524 = n2872 & ~n8523;
  assign n8525 = ~n8520 & n8524;
  assign n8529 = x1136 ^ x876;
  assign n8530 = n8529 ^ x876;
  assign n8531 = x876 ^ x748;
  assign n8532 = n8530 & n8531;
  assign n8533 = n8532 ^ x876;
  assign n8526 = x803 ^ x623;
  assign n8527 = ~x1136 & ~n8526;
  assign n8528 = n8527 ^ x623;
  assign n8534 = n8533 ^ n8528;
  assign n8535 = x1134 & n8534;
  assign n8536 = n8535 ^ n8528;
  assign n8537 = n8536 ^ x1135;
  assign n8538 = n8537 ^ n8536;
  assign n8539 = x789 ^ x710;
  assign n8540 = ~x1136 & n8539;
  assign n8541 = n8540 ^ x710;
  assign n8542 = n8541 ^ x1134;
  assign n8543 = n8542 ^ n8541;
  assign n8544 = n8543 ^ x1135;
  assign n8545 = x1136 ^ x730;
  assign n8546 = x1136 & n8545;
  assign n8547 = n8546 ^ n8541;
  assign n8548 = n8547 ^ x1136;
  assign n8549 = n8544 & n8548;
  assign n8550 = n8549 ^ n8546;
  assign n8551 = n8550 ^ x1136;
  assign n8552 = n8551 ^ n8536;
  assign n8553 = n8538 & n8552;
  assign n8554 = n8553 ^ n8536;
  assign n8555 = n8043 & n8554;
  assign n8556 = ~n8525 & ~n8555;
  assign n8584 = x361 & n8033;
  assign n8585 = x592 ^ x410;
  assign n8586 = n8585 ^ x410;
  assign n8587 = x410 ^ x386;
  assign n8588 = n8586 & n8587;
  assign n8589 = n8588 ^ x410;
  assign n8590 = n7431 & n8589;
  assign n8591 = n3754 & n8590;
  assign n8592 = x434 & n8028;
  assign n8593 = ~n8591 & ~n8592;
  assign n8594 = ~n8584 & n8593;
  assign n8595 = n8594 ^ n1536;
  assign n8596 = n8595 ^ n8594;
  assign n8597 = x199 & n6432;
  assign n8598 = n8597 ^ x293;
  assign n8599 = n8598 ^ n8594;
  assign n8600 = ~n8596 & ~n8599;
  assign n8601 = n8600 ^ n8594;
  assign n8560 = x812 ^ x606;
  assign n8561 = ~x1136 & ~n8560;
  assign n8562 = n8561 ^ x606;
  assign n8557 = x881 ^ x746;
  assign n8558 = ~x1136 & n8557;
  assign n8559 = n8558 ^ x746;
  assign n8563 = n8562 ^ n8559;
  assign n8564 = ~x1134 & n8563;
  assign n8565 = n8564 ^ n8559;
  assign n8566 = n8565 ^ x1135;
  assign n8567 = n8566 ^ n8565;
  assign n8568 = x787 ^ x643;
  assign n8569 = ~x1136 & n8568;
  assign n8570 = n8569 ^ x643;
  assign n8571 = n8570 ^ x1134;
  assign n8572 = n8571 ^ n8570;
  assign n8573 = n8572 ^ x1135;
  assign n8574 = x1136 ^ x729;
  assign n8575 = x1136 & n8574;
  assign n8576 = n8575 ^ n8570;
  assign n8577 = n8576 ^ x1136;
  assign n8578 = n8573 & n8577;
  assign n8579 = n8578 ^ n8575;
  assign n8580 = n8579 ^ x1136;
  assign n8581 = n8580 ^ n8565;
  assign n8582 = n8567 & n8581;
  assign n8583 = n8582 ^ n8565;
  assign n8602 = n8601 ^ n8583;
  assign n8603 = n8602 ^ n8601;
  assign n8604 = n8601 ^ n8042;
  assign n8605 = n8604 ^ n8601;
  assign n8606 = n8603 & n8605;
  assign n8607 = n8606 ^ n8601;
  assign n8608 = ~n2872 & ~n8607;
  assign n8609 = n8608 ^ n8601;
  assign n8610 = x344 & n8033;
  assign n8611 = x592 ^ x366;
  assign n8612 = n8611 ^ x366;
  assign n8613 = x366 ^ x335;
  assign n8614 = ~n8612 & n8613;
  assign n8615 = n8614 ^ x366;
  assign n8616 = n7431 & n8615;
  assign n8617 = n3754 & n8616;
  assign n8618 = x416 & n8028;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = ~n8610 & n8619;
  assign n8621 = n8620 ^ n1536;
  assign n8622 = n8621 ^ n8620;
  assign n8623 = x1069 ^ x259;
  assign n8624 = x199 & n8623;
  assign n8625 = n8624 ^ x259;
  assign n8626 = n8625 ^ n8620;
  assign n8627 = ~n8622 & ~n8626;
  assign n8628 = n8627 ^ n8620;
  assign n8629 = n8628 ^ n8042;
  assign n8630 = n8629 ^ n8628;
  assign n8631 = x870 & n8300;
  assign n8632 = ~x1135 & n4766;
  assign n8633 = n8632 ^ x704;
  assign n8634 = n8633 ^ x1134;
  assign n8635 = n8634 ^ n8633;
  assign n8636 = x635 ^ x620;
  assign n8637 = x1135 & ~n8636;
  assign n8638 = n8637 ^ x620;
  assign n8639 = n8638 ^ n8633;
  assign n8640 = ~n8635 & ~n8639;
  assign n8641 = n8640 ^ n8633;
  assign n8642 = x1136 & ~n8641;
  assign n8643 = ~n8631 & ~n8642;
  assign n8644 = n8643 ^ n8628;
  assign n8645 = n8644 ^ n8628;
  assign n8646 = n8630 & ~n8645;
  assign n8647 = n8646 ^ n8628;
  assign n8648 = ~n2872 & ~n8647;
  assign n8649 = n8648 ^ n8628;
  assign n8654 = x1135 ^ x632;
  assign n8655 = n8654 ^ x632;
  assign n8656 = x632 ^ x613;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = n8657 ^ x632;
  assign n8650 = x1135 ^ x760;
  assign n8651 = n8650 ^ x760;
  assign n8652 = n4799 & n8651;
  assign n8653 = n8652 ^ x760;
  assign n8659 = n8658 ^ n8653;
  assign n8660 = ~x1134 & n8659;
  assign n8661 = n8660 ^ n8653;
  assign n8662 = x1136 & ~n8661;
  assign n8663 = x856 & n8300;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = n8043 & ~n8664;
  assign n8666 = x393 & n2703;
  assign n8667 = x346 & n2806;
  assign n8668 = ~n8666 & ~n8667;
  assign n8669 = x368 & ~x590;
  assign n8670 = ~x591 & n8669;
  assign n8671 = n8668 & ~n8670;
  assign n8672 = n8032 & ~n8671;
  assign n8673 = x418 & n8028;
  assign n8674 = n1536 & ~n8673;
  assign n8675 = ~n8672 & n8674;
  assign n8676 = x1067 ^ x260;
  assign n8677 = x199 & n8676;
  assign n8678 = n8677 ^ x260;
  assign n8679 = ~n1536 & ~n8678;
  assign n8680 = n2872 & ~n8679;
  assign n8681 = ~n8675 & n8680;
  assign n8682 = ~n8665 & ~n8681;
  assign n8683 = x592 ^ x413;
  assign n8684 = n8683 ^ x413;
  assign n8685 = x413 ^ x389;
  assign n8686 = n8684 & n8685;
  assign n8687 = n8686 ^ x413;
  assign n8688 = n7431 & n8687;
  assign n8689 = n3754 & n8688;
  assign n8690 = x438 & n8028;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = n1536 & n8691;
  assign n8693 = x450 & n8033;
  assign n8694 = n8692 & ~n8693;
  assign n8695 = x1036 ^ x255;
  assign n8696 = x199 & n8695;
  assign n8697 = n8696 ^ x255;
  assign n8698 = ~n1536 & ~n8697;
  assign n8699 = n2872 & ~n8698;
  assign n8700 = ~n8694 & n8699;
  assign n8704 = x874 ^ x739;
  assign n8705 = ~x1136 & n8704;
  assign n8706 = n8705 ^ x739;
  assign n8701 = x810 ^ x621;
  assign n8702 = ~x1136 & n8701;
  assign n8703 = n8702 ^ x621;
  assign n8707 = n8706 ^ n8703;
  assign n8708 = x1134 & n8707;
  assign n8709 = n8708 ^ n8703;
  assign n8710 = n8709 ^ x1135;
  assign n8711 = n8710 ^ n8709;
  assign n8712 = x791 ^ x665;
  assign n8713 = ~x1136 & n8712;
  assign n8714 = n8713 ^ x665;
  assign n8715 = n8714 ^ x1134;
  assign n8716 = n8715 ^ n8714;
  assign n8717 = n8716 ^ x1135;
  assign n8718 = x1136 ^ x690;
  assign n8719 = x1136 & n8718;
  assign n8720 = n8719 ^ n8714;
  assign n8721 = n8720 ^ x1136;
  assign n8722 = n8717 & n8721;
  assign n8723 = n8722 ^ n8719;
  assign n8724 = n8723 ^ x1136;
  assign n8725 = n8724 ^ n8709;
  assign n8726 = n8711 & n8725;
  assign n8727 = n8726 ^ n8709;
  assign n8728 = n8043 & n8727;
  assign n8729 = ~n8700 & ~n8728;
  assign n8730 = n7788 ^ x680;
  assign n8731 = n8730 ^ x680;
  assign n8732 = x1100 ^ x680;
  assign n8733 = n8731 & n8732;
  assign n8734 = n8733 ^ x680;
  assign n8735 = ~x962 & n8734;
  assign n8736 = n7788 ^ x681;
  assign n8737 = n8736 ^ x681;
  assign n8738 = x1103 ^ x681;
  assign n8739 = n8737 & n8738;
  assign n8740 = n8739 ^ x681;
  assign n8741 = ~x962 & n8740;
  assign n8742 = x592 ^ x392;
  assign n8743 = n8742 ^ x392;
  assign n8744 = x392 ^ x367;
  assign n8745 = n8743 & n8744;
  assign n8746 = n8745 ^ x392;
  assign n8747 = n7431 & n8746;
  assign n8748 = n3754 & n8747;
  assign n8749 = x417 & n8028;
  assign n8750 = ~n8748 & ~n8749;
  assign n8751 = n1536 & n8750;
  assign n8752 = x345 & n8033;
  assign n8753 = n8751 & ~n8752;
  assign n8754 = x1039 ^ x251;
  assign n8755 = x199 & n8754;
  assign n8756 = n8755 ^ x251;
  assign n8757 = ~n1536 & ~n8756;
  assign n8758 = n2872 & ~n8757;
  assign n8759 = ~n8753 & n8758;
  assign n8764 = x1135 ^ x631;
  assign n8765 = n8764 ^ x631;
  assign n8766 = x631 ^ x610;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = n8767 ^ x631;
  assign n8760 = x1135 ^ x757;
  assign n8761 = n8760 ^ x757;
  assign n8762 = n4777 & n8761;
  assign n8763 = n8762 ^ x757;
  assign n8769 = n8768 ^ n8763;
  assign n8770 = ~x1134 & n8769;
  assign n8771 = n8770 ^ n8763;
  assign n8772 = x1136 & ~n8771;
  assign n8773 = x848 & n8300;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = n8043 & ~n8774;
  assign n8776 = ~n8759 & ~n8775;
  assign n8777 = x953 & n7787;
  assign n8778 = n8777 ^ x684;
  assign n8779 = n8778 ^ x684;
  assign n8780 = x1130 ^ x684;
  assign n8781 = n8779 & ~n8780;
  assign n8782 = n8781 ^ x684;
  assign n8783 = ~x962 & ~n8782;
  assign n8784 = x592 ^ x406;
  assign n8785 = n8784 ^ x406;
  assign n8786 = x406 ^ x382;
  assign n8787 = n8785 & n8786;
  assign n8788 = n8787 ^ x406;
  assign n8789 = n7431 & n8788;
  assign n8790 = n3754 & n8789;
  assign n8791 = x430 & n8028;
  assign n8792 = ~n8790 & ~n8791;
  assign n8793 = n1536 & n8792;
  assign n8794 = x357 & n8033;
  assign n8795 = n8793 & ~n8794;
  assign n8796 = x1076 ^ x199;
  assign n8797 = n8796 ^ x1076;
  assign n8798 = n6142 ^ x1076;
  assign n8799 = ~n8797 & n8798;
  assign n8800 = n8799 ^ x1076;
  assign n8801 = ~n1536 & ~n8800;
  assign n8802 = n2872 & ~n8801;
  assign n8803 = ~n8795 & n8802;
  assign n8814 = x1135 ^ x657;
  assign n8815 = n8814 ^ x657;
  assign n8816 = x657 ^ x652;
  assign n8817 = ~n8815 & ~n8816;
  assign n8818 = n8817 ^ x657;
  assign n8809 = x1135 ^ x744;
  assign n8810 = n8809 ^ x744;
  assign n8811 = x744 ^ x728;
  assign n8812 = n8810 & n8811;
  assign n8813 = n8812 ^ x744;
  assign n8819 = n8818 ^ n8813;
  assign n8820 = ~x1134 & n8819;
  assign n8821 = n8820 ^ n8813;
  assign n8804 = x1134 ^ x860;
  assign n8805 = n8804 ^ x860;
  assign n8806 = x860 ^ x813;
  assign n8807 = ~n8805 & n8806;
  assign n8808 = n8807 ^ x860;
  assign n8822 = n8821 ^ n8808;
  assign n8823 = n8822 ^ n8821;
  assign n8824 = n8821 ^ x1135;
  assign n8825 = n8824 ^ n8821;
  assign n8826 = n8823 & ~n8825;
  assign n8827 = n8826 ^ n8821;
  assign n8828 = ~x1136 & ~n8827;
  assign n8829 = n8828 ^ n8821;
  assign n8830 = n8043 & ~n8829;
  assign n8831 = ~n8803 & ~n8830;
  assign n8832 = n8777 ^ x686;
  assign n8833 = n8832 ^ x686;
  assign n8834 = x1113 ^ x686;
  assign n8835 = n8833 & ~n8834;
  assign n8836 = n8835 ^ x686;
  assign n8837 = ~x962 & ~n8836;
  assign n8838 = n8777 ^ x687;
  assign n8839 = n8838 ^ x687;
  assign n8840 = x1127 ^ x687;
  assign n8841 = n8839 & n8840;
  assign n8842 = n8841 ^ x687;
  assign n8843 = ~x962 & n8842;
  assign n8844 = n8777 ^ x688;
  assign n8845 = n8844 ^ x688;
  assign n8846 = x1115 ^ x688;
  assign n8847 = n8845 & ~n8846;
  assign n8848 = n8847 ^ x688;
  assign n8849 = ~x962 & ~n8848;
  assign n8850 = x351 & n8033;
  assign n8851 = x592 ^ x401;
  assign n8852 = n8851 ^ x401;
  assign n8853 = x401 ^ x376;
  assign n8854 = n8852 & n8853;
  assign n8855 = n8854 ^ x401;
  assign n8856 = n7431 & n8855;
  assign n8857 = n3754 & n8856;
  assign n8858 = x426 & n8028;
  assign n8859 = ~n8857 & ~n8858;
  assign n8860 = ~n8850 & n8859;
  assign n8861 = n8860 ^ n1536;
  assign n8862 = n8861 ^ n8860;
  assign n8863 = x1079 ^ x199;
  assign n8864 = n8863 ^ x1079;
  assign n8865 = n6112 ^ x1079;
  assign n8866 = ~n8864 & n8865;
  assign n8867 = n8866 ^ x1079;
  assign n8868 = n8867 ^ n8860;
  assign n8869 = ~n8862 & ~n8868;
  assign n8870 = n8869 ^ n8860;
  assign n8871 = n8870 ^ n8042;
  assign n8872 = n8871 ^ n8870;
  assign n8881 = x1134 ^ x843;
  assign n8882 = n8881 ^ x843;
  assign n8883 = x843 ^ x798;
  assign n8884 = ~n8882 & n8883;
  assign n8885 = n8884 ^ x843;
  assign n8875 = x658 ^ x655;
  assign n8876 = ~x1135 & ~n8875;
  assign n8877 = n8876 ^ x655;
  assign n8873 = ~x1135 & ~n4872;
  assign n8874 = n8873 ^ x703;
  assign n8878 = n8877 ^ n8874;
  assign n8879 = ~x1134 & ~n8878;
  assign n8880 = n8879 ^ n8874;
  assign n8886 = n8885 ^ n8880;
  assign n8887 = n8886 ^ n8880;
  assign n8888 = n8880 ^ x1135;
  assign n8889 = n8888 ^ n8880;
  assign n8890 = n8887 & ~n8889;
  assign n8891 = n8890 ^ n8880;
  assign n8892 = ~x1136 & n8891;
  assign n8893 = n8892 ^ n8880;
  assign n8894 = n8893 ^ n8870;
  assign n8895 = n8894 ^ n8870;
  assign n8896 = n8872 & n8895;
  assign n8897 = n8896 ^ n8870;
  assign n8898 = ~n2872 & ~n8897;
  assign n8899 = n8898 ^ n8870;
  assign n8900 = n8777 ^ x690;
  assign n8901 = n8900 ^ x690;
  assign n8902 = x1108 ^ x690;
  assign n8903 = n8901 & n8902;
  assign n8904 = n8903 ^ x690;
  assign n8905 = ~x962 & n8904;
  assign n8906 = n8777 ^ x691;
  assign n8907 = n8906 ^ x691;
  assign n8908 = x1107 ^ x691;
  assign n8909 = n8907 & n8908;
  assign n8910 = n8909 ^ x691;
  assign n8911 = ~x962 & n8910;
  assign n8912 = x592 ^ x402;
  assign n8913 = n8912 ^ x402;
  assign n8914 = x402 ^ x317;
  assign n8915 = n8913 & n8914;
  assign n8916 = n8915 ^ x402;
  assign n8917 = n7431 & n8916;
  assign n8918 = n3754 & n8917;
  assign n8919 = x427 & n8028;
  assign n8920 = ~n8918 & ~n8919;
  assign n8921 = n1536 & n8920;
  assign n8922 = x352 & n8033;
  assign n8923 = n8921 & ~n8922;
  assign n8924 = x1078 ^ x199;
  assign n8925 = n8924 ^ x1078;
  assign n8926 = n6124 ^ x1078;
  assign n8927 = ~n8925 & n8926;
  assign n8928 = n8927 ^ x1078;
  assign n8929 = ~n1536 & ~n8928;
  assign n8930 = n2872 & ~n8929;
  assign n8931 = ~n8923 & n8930;
  assign n8940 = x1134 ^ x844;
  assign n8941 = n8940 ^ x844;
  assign n8942 = x844 ^ x801;
  assign n8943 = ~n8941 & n8942;
  assign n8944 = n8943 ^ x844;
  assign n8934 = x656 ^ x649;
  assign n8935 = ~x1135 & ~n8934;
  assign n8936 = n8935 ^ x649;
  assign n8932 = ~x1135 & ~n4682;
  assign n8933 = n8932 ^ x726;
  assign n8937 = n8936 ^ n8933;
  assign n8938 = ~x1134 & ~n8937;
  assign n8939 = n8938 ^ n8933;
  assign n8945 = n8944 ^ n8939;
  assign n8946 = n8945 ^ n8939;
  assign n8947 = n8939 ^ x1135;
  assign n8948 = n8947 ^ n8939;
  assign n8949 = n8946 & ~n8948;
  assign n8950 = n8949 ^ n8939;
  assign n8951 = ~x1136 & n8950;
  assign n8952 = n8951 ^ n8939;
  assign n8953 = n8043 & n8952;
  assign n8954 = ~n8931 & ~n8953;
  assign n8955 = n7788 ^ x693;
  assign n8956 = n8955 ^ x693;
  assign n8957 = x1129 ^ x693;
  assign n8958 = n8956 & ~n8957;
  assign n8959 = n8958 ^ x693;
  assign n8960 = ~x962 & ~n8959;
  assign n8961 = n8777 ^ x694;
  assign n8962 = n8961 ^ x694;
  assign n8963 = x1128 ^ x694;
  assign n8964 = n8962 & ~n8963;
  assign n8965 = n8964 ^ x694;
  assign n8966 = ~x962 & ~n8965;
  assign n8967 = n7788 ^ x695;
  assign n8968 = n8967 ^ x695;
  assign n8969 = x1111 ^ x695;
  assign n8970 = n8968 & ~n8969;
  assign n8971 = n8970 ^ x695;
  assign n8972 = ~x962 & ~n8971;
  assign n8973 = n8777 ^ x696;
  assign n8974 = n8973 ^ x696;
  assign n8975 = x1100 ^ x696;
  assign n8976 = n8974 & n8975;
  assign n8977 = n8976 ^ x696;
  assign n8978 = ~x962 & n8977;
  assign n8979 = n8777 ^ x697;
  assign n8980 = n8979 ^ x697;
  assign n8981 = x1129 ^ x697;
  assign n8982 = n8980 & ~n8981;
  assign n8983 = n8982 ^ x697;
  assign n8984 = ~x962 & ~n8983;
  assign n8985 = n8777 ^ x698;
  assign n8986 = n8985 ^ x698;
  assign n8987 = x1116 ^ x698;
  assign n8988 = n8986 & ~n8987;
  assign n8989 = n8988 ^ x698;
  assign n8990 = ~x962 & ~n8989;
  assign n8991 = n8777 ^ x699;
  assign n8992 = n8991 ^ x699;
  assign n8993 = x1103 ^ x699;
  assign n8994 = n8992 & n8993;
  assign n8995 = n8994 ^ x699;
  assign n8996 = ~x962 & n8995;
  assign n8997 = n8777 ^ x700;
  assign n8998 = n8997 ^ x700;
  assign n8999 = x1110 ^ x700;
  assign n9000 = n8998 & n8999;
  assign n9001 = n9000 ^ x700;
  assign n9002 = ~x962 & n9001;
  assign n9003 = n8777 ^ x701;
  assign n9004 = n9003 ^ x701;
  assign n9005 = x1123 ^ x701;
  assign n9006 = n9004 & ~n9005;
  assign n9007 = n9006 ^ x701;
  assign n9008 = ~x962 & ~n9007;
  assign n9009 = n8777 ^ x702;
  assign n9010 = n9009 ^ x702;
  assign n9011 = x1117 ^ x702;
  assign n9012 = n9010 & ~n9011;
  assign n9013 = n9012 ^ x702;
  assign n9014 = ~x962 & ~n9013;
  assign n9015 = n8777 ^ x703;
  assign n9016 = n9015 ^ x703;
  assign n9017 = x1124 ^ x703;
  assign n9018 = n9016 & n9017;
  assign n9019 = n9018 ^ x703;
  assign n9020 = ~x962 & n9019;
  assign n9021 = n8777 ^ x704;
  assign n9022 = n9021 ^ x704;
  assign n9023 = x1112 ^ x704;
  assign n9024 = n9022 & ~n9023;
  assign n9025 = n9024 ^ x704;
  assign n9026 = ~x962 & ~n9025;
  assign n9027 = n8777 ^ x705;
  assign n9028 = n9027 ^ x705;
  assign n9029 = x1125 ^ x705;
  assign n9030 = n9028 & n9029;
  assign n9031 = n9030 ^ x705;
  assign n9032 = ~x962 & n9031;
  assign n9033 = n8777 ^ x706;
  assign n9034 = n9033 ^ x706;
  assign n9035 = x1105 ^ x706;
  assign n9036 = n9034 & n9035;
  assign n9037 = n9036 ^ x706;
  assign n9038 = ~x962 & n9037;
  assign n9039 = x592 ^ x395;
  assign n9040 = n9039 ^ x395;
  assign n9041 = x395 ^ x370;
  assign n9042 = n9040 & n9041;
  assign n9043 = n9042 ^ x395;
  assign n9044 = n7431 & n9043;
  assign n9045 = n3754 & n9044;
  assign n9046 = x420 & n8028;
  assign n9047 = ~n9045 & ~n9046;
  assign n9048 = n1536 & n9047;
  assign n9049 = x347 & n8033;
  assign n9050 = n9048 & ~n9049;
  assign n9052 = x1055 ^ x1048;
  assign n9051 = x1055 ^ x304;
  assign n9053 = n9052 ^ n9051;
  assign n9054 = n9051 ^ x200;
  assign n9055 = n9054 ^ n9051;
  assign n9056 = n9053 & n9055;
  assign n9057 = n9056 ^ n9051;
  assign n9058 = ~x199 & n9057;
  assign n9059 = n9058 ^ x1055;
  assign n9060 = ~n1536 & ~n9059;
  assign n9061 = n2872 & ~n9060;
  assign n9062 = ~n9050 & n9061;
  assign n9063 = x847 & n8300;
  assign n9064 = ~x1135 & n4810;
  assign n9065 = n9064 ^ x702;
  assign n9066 = n9065 ^ x1134;
  assign n9067 = n9066 ^ n9065;
  assign n9068 = x627 ^ x618;
  assign n9069 = x1135 & n9068;
  assign n9070 = n9069 ^ x618;
  assign n9071 = n9070 ^ n9065;
  assign n9072 = ~n9067 & ~n9071;
  assign n9073 = n9072 ^ n9065;
  assign n9074 = x1136 & ~n9073;
  assign n9075 = ~n9063 & ~n9074;
  assign n9076 = n8043 & ~n9075;
  assign n9077 = ~n9062 & ~n9076;
  assign n9078 = x321 & n8033;
  assign n9079 = x592 ^ x442;
  assign n9080 = n9079 ^ x442;
  assign n9081 = x442 ^ x328;
  assign n9082 = ~n9080 & n9081;
  assign n9083 = n9082 ^ x442;
  assign n9084 = n7431 & n9083;
  assign n9085 = n3754 & n9084;
  assign n9086 = x459 & n8028;
  assign n9087 = ~n9085 & ~n9086;
  assign n9088 = ~n9078 & n9087;
  assign n9089 = n9088 ^ n1536;
  assign n9090 = n9089 ^ n9088;
  assign n9092 = x1084 ^ x1058;
  assign n9091 = x1058 ^ x305;
  assign n9093 = n9092 ^ n9091;
  assign n9094 = n9091 ^ x200;
  assign n9095 = n9094 ^ n9091;
  assign n9096 = n9093 & n9095;
  assign n9097 = n9096 ^ n9091;
  assign n9098 = ~x199 & n9097;
  assign n9099 = n9098 ^ x1058;
  assign n9100 = n9099 ^ n9088;
  assign n9101 = ~n9090 & ~n9100;
  assign n9102 = n9101 ^ n9088;
  assign n9103 = n9102 ^ n8042;
  assign n9104 = n9103 ^ n9102;
  assign n9105 = x857 & n8300;
  assign n9106 = ~x1135 & n4821;
  assign n9107 = n9106 ^ x709;
  assign n9108 = n9107 ^ x1134;
  assign n9109 = n9108 ^ n9107;
  assign n9110 = x660 ^ x609;
  assign n9111 = x1135 & n9110;
  assign n9112 = n9111 ^ x609;
  assign n9113 = n9112 ^ n9107;
  assign n9114 = ~n9109 & ~n9113;
  assign n9115 = n9114 ^ n9107;
  assign n9116 = x1136 & ~n9115;
  assign n9117 = ~n9105 & ~n9116;
  assign n9118 = n9117 ^ n9102;
  assign n9119 = n9118 ^ n9102;
  assign n9120 = n9104 & ~n9119;
  assign n9121 = n9120 ^ n9102;
  assign n9122 = ~n2872 & ~n9121;
  assign n9123 = n9122 ^ n9102;
  assign n9124 = n8777 ^ x709;
  assign n9125 = n9124 ^ x709;
  assign n9126 = x1118 ^ x709;
  assign n9127 = n9125 & ~n9126;
  assign n9128 = n9127 ^ x709;
  assign n9129 = ~x962 & ~n9128;
  assign n9130 = n7788 ^ x710;
  assign n9131 = n9130 ^ x710;
  assign n9132 = x1106 ^ x710;
  assign n9133 = n9131 & n9132;
  assign n9134 = n9133 ^ x710;
  assign n9135 = ~x962 & n9134;
  assign n9136 = x592 ^ x398;
  assign n9137 = n9136 ^ x398;
  assign n9138 = x398 ^ x373;
  assign n9139 = n9137 & n9138;
  assign n9140 = n9139 ^ x398;
  assign n9141 = n7431 & n9140;
  assign n9142 = n3754 & n9141;
  assign n9143 = x423 & n8028;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = n1536 & n9144;
  assign n9146 = x348 & n8033;
  assign n9147 = n9145 & ~n9146;
  assign n9149 = x1087 ^ x306;
  assign n9148 = x1087 ^ x1059;
  assign n9150 = n9149 ^ n9148;
  assign n9151 = n9149 ^ x200;
  assign n9152 = n9151 ^ n9149;
  assign n9153 = n9150 & n9152;
  assign n9154 = n9153 ^ n9149;
  assign n9155 = ~x199 & n9154;
  assign n9156 = n9155 ^ x1087;
  assign n9157 = ~n1536 & ~n9156;
  assign n9158 = n2872 & ~n9157;
  assign n9159 = ~n9147 & n9158;
  assign n9160 = x858 & n8300;
  assign n9161 = ~x1135 & n4711;
  assign n9162 = n9161 ^ x725;
  assign n9163 = n9162 ^ x1134;
  assign n9164 = n9163 ^ n9162;
  assign n9165 = x647 ^ x630;
  assign n9166 = x1135 & n9165;
  assign n9167 = n9166 ^ x630;
  assign n9168 = n9167 ^ n9162;
  assign n9169 = ~n9164 & ~n9168;
  assign n9170 = n9169 ^ n9162;
  assign n9171 = x1136 & ~n9170;
  assign n9172 = ~n9160 & ~n9171;
  assign n9173 = n8043 & ~n9172;
  assign n9174 = ~n9159 & ~n9173;
  assign n9175 = x592 ^ x400;
  assign n9176 = n9175 ^ x400;
  assign n9177 = x400 ^ x374;
  assign n9178 = n9176 & n9177;
  assign n9179 = n9178 ^ x400;
  assign n9180 = n7431 & n9179;
  assign n9181 = n3754 & n9180;
  assign n9182 = x425 & n8028;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = n1536 & n9183;
  assign n9185 = x350 & n8033;
  assign n9186 = n9184 & ~n9185;
  assign n9188 = x1044 ^ x1035;
  assign n9187 = x1035 ^ x298;
  assign n9189 = n9188 ^ n9187;
  assign n9190 = n9187 ^ x200;
  assign n9191 = n9190 ^ n9187;
  assign n9192 = n9189 & n9191;
  assign n9193 = n9192 ^ n9187;
  assign n9194 = ~x199 & n9193;
  assign n9195 = n9194 ^ x1035;
  assign n9196 = ~n1536 & ~n9195;
  assign n9197 = n2872 & ~n9196;
  assign n9198 = ~n9186 & n9197;
  assign n9199 = x842 & n8300;
  assign n9200 = ~x1135 & n4722;
  assign n9201 = n9200 ^ x701;
  assign n9202 = n9201 ^ x1134;
  assign n9203 = n9202 ^ n9201;
  assign n9204 = x715 ^ x644;
  assign n9205 = x1135 & n9204;
  assign n9206 = n9205 ^ x644;
  assign n9207 = n9206 ^ n9201;
  assign n9208 = ~n9203 & ~n9207;
  assign n9209 = n9208 ^ n9201;
  assign n9210 = x1136 & ~n9209;
  assign n9211 = ~n9199 & ~n9210;
  assign n9212 = n8043 & ~n9211;
  assign n9213 = ~n9198 & ~n9212;
  assign n9214 = x592 ^ x396;
  assign n9215 = n9214 ^ x396;
  assign n9216 = x396 ^ x371;
  assign n9217 = n9215 & n9216;
  assign n9218 = n9217 ^ x396;
  assign n9219 = n7431 & n9218;
  assign n9220 = n3754 & n9219;
  assign n9221 = x421 & n8028;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = n1536 & n9222;
  assign n9224 = x322 & n8033;
  assign n9225 = n9223 & ~n9224;
  assign n9227 = x1051 ^ x309;
  assign n9226 = x1072 ^ x1051;
  assign n9228 = n9227 ^ n9226;
  assign n9229 = n9227 ^ x200;
  assign n9230 = n9229 ^ n9227;
  assign n9231 = n9228 & n9230;
  assign n9232 = n9231 ^ n9227;
  assign n9233 = ~x199 & n9232;
  assign n9234 = n9233 ^ x1051;
  assign n9235 = ~n1536 & ~n9234;
  assign n9236 = n2872 & ~n9235;
  assign n9237 = ~n9225 & n9236;
  assign n9238 = x854 & n8300;
  assign n9239 = ~x1135 & n4832;
  assign n9240 = n9239 ^ x734;
  assign n9241 = n9240 ^ x1134;
  assign n9242 = n9241 ^ n9240;
  assign n9243 = x629 ^ x628;
  assign n9244 = ~x1135 & n9243;
  assign n9245 = n9244 ^ x628;
  assign n9246 = n9245 ^ n9240;
  assign n9247 = ~n9242 & ~n9246;
  assign n9248 = n9247 ^ n9240;
  assign n9249 = x1136 & ~n9248;
  assign n9250 = ~n9238 & ~n9249;
  assign n9251 = n8043 & ~n9250;
  assign n9252 = ~n9237 & ~n9251;
  assign n9253 = x461 & n8033;
  assign n9254 = x592 ^ x439;
  assign n9255 = n9254 ^ x439;
  assign n9256 = x439 ^ x326;
  assign n9257 = ~n9255 & n9256;
  assign n9258 = n9257 ^ x439;
  assign n9259 = n7431 & n9258;
  assign n9260 = n3754 & n9259;
  assign n9261 = x449 & n8028;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~n9253 & n9262;
  assign n9264 = n9263 ^ n1536;
  assign n9265 = n9264 ^ n9263;
  assign n9266 = x1057 ^ x199;
  assign n9267 = n9266 ^ x1057;
  assign n9268 = n6076 ^ x1057;
  assign n9269 = ~n9267 & n9268;
  assign n9270 = n9269 ^ x1057;
  assign n9271 = n9270 ^ n9263;
  assign n9272 = ~n9265 & ~n9271;
  assign n9273 = n9272 ^ n9263;
  assign n9274 = n9273 ^ n8042;
  assign n9275 = n9274 ^ n9273;
  assign n9286 = x1135 ^ x693;
  assign n9287 = n9286 ^ x693;
  assign n9288 = x693 ^ x653;
  assign n9289 = ~n9287 & ~n9288;
  assign n9290 = n9289 ^ x693;
  assign n9281 = x1135 ^ x762;
  assign n9282 = n9281 ^ x762;
  assign n9283 = x762 ^ x697;
  assign n9284 = n9282 & n9283;
  assign n9285 = n9284 ^ x762;
  assign n9291 = n9290 ^ n9285;
  assign n9292 = ~x1134 & n9291;
  assign n9293 = n9292 ^ n9285;
  assign n9276 = x1134 ^ x867;
  assign n9277 = n9276 ^ x867;
  assign n9278 = x867 ^ x816;
  assign n9279 = ~n9277 & n9278;
  assign n9280 = n9279 ^ x867;
  assign n9294 = n9293 ^ n9280;
  assign n9295 = n9294 ^ n9293;
  assign n9296 = n9293 ^ x1135;
  assign n9297 = n9296 ^ n9293;
  assign n9298 = n9295 & ~n9297;
  assign n9299 = n9298 ^ n9293;
  assign n9300 = ~x1136 & ~n9299;
  assign n9301 = n9300 ^ n9293;
  assign n9302 = n9301 ^ n9273;
  assign n9303 = n9302 ^ n9273;
  assign n9304 = n9275 & ~n9303;
  assign n9305 = n9304 ^ n9273;
  assign n9306 = ~n2872 & ~n9305;
  assign n9307 = n9306 ^ n9273;
  assign n9308 = n7788 ^ x715;
  assign n9309 = n9308 ^ x715;
  assign n9310 = x1123 ^ x715;
  assign n9311 = n9309 & n9310;
  assign n9312 = n9311 ^ x715;
  assign n9313 = ~x962 & n9312;
  assign n9314 = x349 & n8033;
  assign n9315 = x592 ^ x440;
  assign n9316 = n9315 ^ x440;
  assign n9317 = x440 ^ x329;
  assign n9318 = ~n9316 & n9317;
  assign n9319 = n9318 ^ x440;
  assign n9320 = n7431 & n9319;
  assign n9321 = n3754 & n9320;
  assign n9322 = ~n9314 & ~n9321;
  assign n9323 = x454 & n8028;
  assign n9324 = n1536 & ~n9323;
  assign n9325 = n9322 & n9324;
  assign n9327 = x1053 ^ x1043;
  assign n9326 = x1043 ^ x307;
  assign n9328 = n9327 ^ n9326;
  assign n9329 = n9326 ^ x200;
  assign n9330 = n9329 ^ n9326;
  assign n9331 = n9328 & n9330;
  assign n9332 = n9331 ^ n9326;
  assign n9333 = ~x199 & n9332;
  assign n9334 = n9333 ^ x1043;
  assign n9335 = ~n1536 & ~n9334;
  assign n9336 = n2872 & ~n9335;
  assign n9337 = ~n9325 & n9336;
  assign n9338 = x845 & n8300;
  assign n9339 = ~x1135 & n4609;
  assign n9340 = n9339 ^ x738;
  assign n9341 = n9340 ^ x1134;
  assign n9342 = n9341 ^ n9340;
  assign n9343 = x641 ^ x626;
  assign n9344 = x1135 & n9343;
  assign n9345 = n9344 ^ x626;
  assign n9346 = n9345 ^ n9340;
  assign n9347 = ~n9342 & ~n9346;
  assign n9348 = n9347 ^ n9340;
  assign n9349 = x1136 & ~n9348;
  assign n9350 = ~n9338 & ~n9349;
  assign n9351 = n8043 & ~n9350;
  assign n9352 = ~n9337 & ~n9351;
  assign n9353 = x462 & n8033;
  assign n9354 = x592 ^ x377;
  assign n9355 = n9354 ^ x377;
  assign n9356 = x377 ^ x318;
  assign n9357 = ~n9355 & n9356;
  assign n9358 = n9357 ^ x377;
  assign n9359 = n7431 & n9358;
  assign n9360 = n3754 & n9359;
  assign n9361 = x448 & n8028;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = ~n9353 & n9362;
  assign n9364 = n9363 ^ n1536;
  assign n9365 = n9364 ^ n9363;
  assign n9366 = x1074 ^ x199;
  assign n9367 = n9366 ^ x1074;
  assign n9368 = n6118 ^ x1074;
  assign n9369 = ~n9367 & n9368;
  assign n9370 = n9369 ^ x1074;
  assign n9371 = n9370 ^ n9363;
  assign n9372 = ~n9365 & ~n9371;
  assign n9373 = n9372 ^ n9363;
  assign n9374 = n9373 ^ n8042;
  assign n9375 = n9374 ^ n9373;
  assign n9386 = x1134 ^ x839;
  assign n9387 = n9386 ^ x839;
  assign n9388 = x839 ^ x800;
  assign n9389 = ~n9387 & n9388;
  assign n9390 = n9389 ^ x839;
  assign n9376 = ~x1135 & ~n4903;
  assign n9377 = n9376 ^ x705;
  assign n9378 = n9377 ^ x1134;
  assign n9379 = n9378 ^ n9377;
  assign n9380 = x669 ^ x645;
  assign n9381 = x1135 & ~n9380;
  assign n9382 = n9381 ^ x645;
  assign n9383 = n9382 ^ n9377;
  assign n9384 = ~n9379 & n9383;
  assign n9385 = n9384 ^ n9377;
  assign n9391 = n9390 ^ n9385;
  assign n9392 = n9391 ^ n9385;
  assign n9393 = n9385 ^ x1135;
  assign n9394 = n9393 ^ n9385;
  assign n9395 = n9392 & ~n9394;
  assign n9396 = n9395 ^ n9385;
  assign n9397 = ~x1136 & n9396;
  assign n9398 = n9397 ^ n9385;
  assign n9399 = n9398 ^ n9373;
  assign n9400 = n9399 ^ n9373;
  assign n9401 = n9375 & n9400;
  assign n9402 = n9401 ^ n9373;
  assign n9403 = ~n2872 & ~n9402;
  assign n9404 = n9403 ^ n9373;
  assign n9405 = x315 & n8033;
  assign n9406 = x419 & n8028;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = x592 ^ x394;
  assign n9409 = n9408 ^ x394;
  assign n9410 = x394 ^ x369;
  assign n9411 = n9409 & n9410;
  assign n9412 = n9411 ^ x394;
  assign n9413 = n7431 & n9412;
  assign n9414 = n3754 & n9413;
  assign n9415 = n1536 & ~n9414;
  assign n9416 = n9407 & n9415;
  assign n9418 = x1080 ^ x303;
  assign n9417 = x1080 ^ x1049;
  assign n9419 = n9418 ^ n9417;
  assign n9420 = n9418 ^ x200;
  assign n9421 = n9420 ^ n9418;
  assign n9422 = n9419 & n9421;
  assign n9423 = n9422 ^ n9418;
  assign n9424 = ~x199 & n9423;
  assign n9425 = n9424 ^ x1080;
  assign n9426 = ~n1536 & ~n9425;
  assign n9427 = n2872 & ~n9426;
  assign n9428 = ~n9416 & n9427;
  assign n9429 = x853 & n8300;
  assign n9430 = ~x1135 & n4664;
  assign n9431 = n9430 ^ x698;
  assign n9432 = n9431 ^ x1134;
  assign n9433 = n9432 ^ n9431;
  assign n9434 = x625 ^ x608;
  assign n9435 = x1135 & n9434;
  assign n9436 = n9435 ^ x608;
  assign n9437 = n9436 ^ n9431;
  assign n9438 = ~n9433 & ~n9437;
  assign n9439 = n9438 ^ n9431;
  assign n9440 = x1136 & ~n9439;
  assign n9441 = ~n9429 & ~n9440;
  assign n9442 = n8043 & ~n9441;
  assign n9443 = ~n9428 & ~n9442;
  assign n9444 = x353 & n8033;
  assign n9445 = x592 ^ x378;
  assign n9446 = n9445 ^ x378;
  assign n9447 = x378 ^ x325;
  assign n9448 = ~n9446 & n9447;
  assign n9449 = n9448 ^ x378;
  assign n9450 = n7431 & n9449;
  assign n9451 = n3754 & n9450;
  assign n9452 = x451 & n8028;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = ~n9444 & n9453;
  assign n9455 = n9454 ^ n1536;
  assign n9456 = n9455 ^ n9454;
  assign n9457 = x1063 ^ x199;
  assign n9458 = n9457 ^ x1063;
  assign n9459 = n6130 ^ x1063;
  assign n9460 = ~n9458 & n9459;
  assign n9461 = n9460 ^ x1063;
  assign n9462 = n9461 ^ n9454;
  assign n9463 = ~n9456 & ~n9462;
  assign n9464 = n9463 ^ n9454;
  assign n9465 = n9464 ^ n8042;
  assign n9466 = n9465 ^ n9464;
  assign n9476 = x1135 ^ x650;
  assign n9477 = n9476 ^ x650;
  assign n9478 = x650 ^ x636;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = n9479 ^ x650;
  assign n9472 = x1135 ^ x774;
  assign n9473 = n9472 ^ x774;
  assign n9474 = ~n4642 & n9473;
  assign n9475 = n9474 ^ x774;
  assign n9481 = n9480 ^ n9475;
  assign n9482 = ~x1134 & n9481;
  assign n9483 = n9482 ^ n9475;
  assign n9467 = x1134 ^ x868;
  assign n9468 = n9467 ^ x868;
  assign n9469 = x868 ^ x807;
  assign n9470 = ~n9468 & n9469;
  assign n9471 = n9470 ^ x868;
  assign n9484 = n9483 ^ n9471;
  assign n9485 = n9484 ^ n9483;
  assign n9486 = n9483 ^ x1135;
  assign n9487 = n9486 ^ n9483;
  assign n9488 = n9485 & ~n9487;
  assign n9489 = n9488 ^ n9483;
  assign n9490 = ~x1136 & ~n9489;
  assign n9491 = n9490 ^ n9483;
  assign n9492 = n9491 ^ n9464;
  assign n9493 = n9492 ^ n9464;
  assign n9494 = n9466 & ~n9493;
  assign n9495 = n9494 ^ n9464;
  assign n9496 = ~n2872 & ~n9495;
  assign n9497 = n9496 ^ n9464;
  assign n9498 = x356 & n8033;
  assign n9499 = x592 ^ x405;
  assign n9500 = n9499 ^ x405;
  assign n9501 = x405 ^ x381;
  assign n9502 = n9500 & n9501;
  assign n9503 = n9502 ^ x405;
  assign n9504 = n7431 & n9503;
  assign n9505 = n3754 & n9504;
  assign n9506 = x445 & n8028;
  assign n9507 = ~n9505 & ~n9506;
  assign n9508 = ~n9498 & n9507;
  assign n9509 = n9508 ^ n1536;
  assign n9510 = n9509 ^ n9508;
  assign n9511 = x1081 ^ x199;
  assign n9512 = n9511 ^ x1081;
  assign n9513 = n6148 ^ x1081;
  assign n9514 = ~n9512 & n9513;
  assign n9515 = n9514 ^ x1081;
  assign n9516 = n9515 ^ n9508;
  assign n9517 = ~n9510 & ~n9516;
  assign n9518 = n9517 ^ n9508;
  assign n9519 = n9518 ^ n8042;
  assign n9520 = n9519 ^ n9518;
  assign n9534 = x1134 ^ x880;
  assign n9535 = n9534 ^ x880;
  assign n9536 = x880 ^ x794;
  assign n9537 = ~n9535 & n9536;
  assign n9538 = n9537 ^ x880;
  assign n9526 = x1135 ^ x654;
  assign n9527 = n9526 ^ x654;
  assign n9528 = x654 ^ x651;
  assign n9529 = ~n9527 & ~n9528;
  assign n9530 = n9529 ^ x654;
  assign n9521 = x1135 ^ x750;
  assign n9522 = n9521 ^ x750;
  assign n9523 = x750 ^ x684;
  assign n9524 = n9522 & n9523;
  assign n9525 = n9524 ^ x750;
  assign n9531 = n9530 ^ n9525;
  assign n9532 = ~x1134 & n9531;
  assign n9533 = n9532 ^ n9525;
  assign n9539 = n9538 ^ n9533;
  assign n9540 = n9539 ^ n9533;
  assign n9541 = n9533 ^ x1135;
  assign n9542 = n9541 ^ n9533;
  assign n9543 = n9540 & ~n9542;
  assign n9544 = n9543 ^ n9533;
  assign n9545 = ~x1136 & ~n9544;
  assign n9546 = n9545 ^ n9533;
  assign n9547 = n9546 ^ n9518;
  assign n9548 = n9547 ^ n9518;
  assign n9549 = n9520 & ~n9548;
  assign n9550 = n9549 ^ n9518;
  assign n9551 = ~n2872 & ~n9550;
  assign n9552 = n9551 ^ n9518;
  assign n9553 = x747 & x773;
  assign n9554 = x731 & ~x945;
  assign n9555 = n9553 & n9554;
  assign n9556 = x775 & x988;
  assign n9557 = n9555 & n9556;
  assign n9558 = x769 & n9557;
  assign n9559 = n9558 ^ x721;
  assign n9560 = x798 ^ x765;
  assign n9561 = x800 ^ x771;
  assign n9562 = ~n9560 & ~n9561;
  assign n9563 = x807 ^ x747;
  assign n9564 = x816 ^ x775;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = n9562 & n9565;
  assign n9567 = x794 ^ x769;
  assign n9568 = x801 ^ x773;
  assign n9569 = ~n9567 & ~n9568;
  assign n9570 = x813 ^ x721;
  assign n9571 = x795 ^ x731;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = n9569 & n9572;
  assign n9574 = n9566 & n9573;
  assign n9575 = n9559 & ~n9574;
  assign n9576 = x592 ^ x403;
  assign n9577 = n9576 ^ x403;
  assign n9578 = x403 ^ x379;
  assign n9579 = n9577 & n9578;
  assign n9580 = n9579 ^ x403;
  assign n9581 = n7431 & n9580;
  assign n9582 = n3754 & n9581;
  assign n9583 = x428 & n8028;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = n1536 & n9584;
  assign n9586 = x354 & n8033;
  assign n9587 = n9585 & ~n9586;
  assign n9588 = x1045 ^ x199;
  assign n9589 = n9588 ^ x1045;
  assign n9590 = n6136 ^ x1045;
  assign n9591 = ~n9589 & n9590;
  assign n9592 = n9591 ^ x1045;
  assign n9593 = ~n1536 & ~n9592;
  assign n9594 = n2872 & ~n9593;
  assign n9595 = ~n9587 & n9594;
  assign n9606 = x1135 ^ x732;
  assign n9607 = n9606 ^ x732;
  assign n9608 = x732 ^ x640;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = n9609 ^ x732;
  assign n9601 = x1135 ^ x776;
  assign n9602 = n9601 ^ x776;
  assign n9603 = x776 ^ x694;
  assign n9604 = n9602 & n9603;
  assign n9605 = n9604 ^ x776;
  assign n9611 = n9610 ^ n9605;
  assign n9612 = ~x1134 & n9611;
  assign n9613 = n9612 ^ n9605;
  assign n9596 = x1134 ^ x851;
  assign n9597 = n9596 ^ x851;
  assign n9598 = x851 ^ x795;
  assign n9599 = ~n9597 & n9598;
  assign n9600 = n9599 ^ x851;
  assign n9614 = n9613 ^ n9600;
  assign n9615 = n9614 ^ n9613;
  assign n9616 = n9613 ^ x1135;
  assign n9617 = n9616 ^ n9613;
  assign n9618 = n9615 & ~n9617;
  assign n9619 = n9618 ^ n9613;
  assign n9620 = ~x1136 & ~n9619;
  assign n9621 = n9620 ^ n9613;
  assign n9622 = n8043 & ~n9621;
  assign n9623 = ~n9595 & ~n9622;
  assign n9624 = n8777 ^ x723;
  assign n9625 = n9624 ^ x723;
  assign n9626 = x1111 ^ x723;
  assign n9627 = n9625 & ~n9626;
  assign n9628 = n9627 ^ x723;
  assign n9629 = ~x962 & ~n9628;
  assign n9630 = n8777 ^ x724;
  assign n9631 = n9630 ^ x724;
  assign n9632 = x1114 ^ x724;
  assign n9633 = n9631 & ~n9632;
  assign n9634 = n9633 ^ x724;
  assign n9635 = ~x962 & ~n9634;
  assign n9636 = n8777 ^ x725;
  assign n9637 = n9636 ^ x725;
  assign n9638 = x1120 ^ x725;
  assign n9639 = n9637 & ~n9638;
  assign n9640 = n9639 ^ x725;
  assign n9641 = ~x962 & ~n9640;
  assign n9642 = n8777 ^ x726;
  assign n9643 = n9642 ^ x726;
  assign n9644 = x1126 ^ x726;
  assign n9645 = n9643 & n9644;
  assign n9646 = n9645 ^ x726;
  assign n9647 = ~x962 & n9646;
  assign n9648 = n8777 ^ x727;
  assign n9649 = n9648 ^ x727;
  assign n9650 = x1102 ^ x727;
  assign n9651 = n9649 & n9650;
  assign n9652 = n9651 ^ x727;
  assign n9653 = ~x962 & n9652;
  assign n9654 = n8777 ^ x728;
  assign n9655 = n9654 ^ x728;
  assign n9656 = x1131 ^ x728;
  assign n9657 = n9655 & ~n9656;
  assign n9658 = n9657 ^ x728;
  assign n9659 = ~x962 & ~n9658;
  assign n9660 = n8777 ^ x729;
  assign n9661 = n9660 ^ x729;
  assign n9662 = x1104 ^ x729;
  assign n9663 = n9661 & n9662;
  assign n9664 = n9663 ^ x729;
  assign n9665 = ~x962 & n9664;
  assign n9666 = n8777 ^ x730;
  assign n9667 = n9666 ^ x730;
  assign n9668 = x1106 ^ x730;
  assign n9669 = n9667 & n9668;
  assign n9670 = n9669 ^ x730;
  assign n9671 = ~x962 & n9670;
  assign n9672 = ~x945 & x988;
  assign n9673 = n9553 & n9672;
  assign n9674 = n9673 ^ x731;
  assign n9675 = ~n9574 & n9674;
  assign n9676 = n7788 ^ x732;
  assign n9677 = n9676 ^ x732;
  assign n9678 = x1128 ^ x732;
  assign n9679 = n9677 & ~n9678;
  assign n9680 = n9679 ^ x732;
  assign n9681 = ~x962 & ~n9680;
  assign n9682 = x316 & n8033;
  assign n9683 = x592 ^ x399;
  assign n9684 = n9683 ^ x399;
  assign n9685 = x399 ^ x375;
  assign n9686 = n9684 & n9685;
  assign n9687 = n9686 ^ x399;
  assign n9688 = n7431 & n9687;
  assign n9689 = n3754 & n9688;
  assign n9690 = x424 & n8028;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = ~n9682 & n9691;
  assign n9693 = n9692 ^ n1536;
  assign n9694 = n9693 ^ n9692;
  assign n9696 = x1047 ^ x1037;
  assign n9695 = x1047 ^ x308;
  assign n9697 = n9696 ^ n9695;
  assign n9698 = n9695 ^ x200;
  assign n9699 = n9698 ^ n9695;
  assign n9700 = n9697 & n9699;
  assign n9701 = n9700 ^ n9695;
  assign n9702 = ~x199 & n9701;
  assign n9703 = n9702 ^ x1047;
  assign n9704 = n9703 ^ n9692;
  assign n9705 = ~n9694 & ~n9704;
  assign n9706 = n9705 ^ n9692;
  assign n9707 = n9706 ^ n8042;
  assign n9708 = n9707 ^ n9706;
  assign n9709 = x838 & n8300;
  assign n9710 = ~x1135 & n4861;
  assign n9711 = n9710 ^ x737;
  assign n9712 = n9711 ^ x1134;
  assign n9713 = n9712 ^ n9711;
  assign n9714 = x648 ^ x619;
  assign n9715 = x1135 & n9714;
  assign n9716 = n9715 ^ x619;
  assign n9717 = n9716 ^ n9711;
  assign n9718 = ~n9713 & ~n9717;
  assign n9719 = n9718 ^ n9711;
  assign n9720 = x1136 & ~n9719;
  assign n9721 = ~n9709 & ~n9720;
  assign n9722 = n9721 ^ n9706;
  assign n9723 = n9722 ^ n9706;
  assign n9724 = n9708 & ~n9723;
  assign n9725 = n9724 ^ n9706;
  assign n9726 = ~n2872 & ~n9725;
  assign n9727 = n9726 ^ n9706;
  assign n9728 = n8777 ^ x734;
  assign n9729 = n9728 ^ x734;
  assign n9730 = x1119 ^ x734;
  assign n9731 = n9729 & ~n9730;
  assign n9732 = n9731 ^ x734;
  assign n9733 = ~x962 & ~n9732;
  assign n9734 = n8777 ^ x735;
  assign n9735 = n9734 ^ x735;
  assign n9736 = x1109 ^ x735;
  assign n9737 = n9735 & n9736;
  assign n9738 = n9737 ^ x735;
  assign n9739 = ~x962 & n9738;
  assign n9740 = n8777 ^ x736;
  assign n9741 = n9740 ^ x736;
  assign n9742 = x1101 ^ x736;
  assign n9743 = n9741 & n9742;
  assign n9744 = n9743 ^ x736;
  assign n9745 = ~x962 & n9744;
  assign n9746 = n8777 ^ x737;
  assign n9747 = n9746 ^ x737;
  assign n9748 = x1122 ^ x737;
  assign n9749 = n9747 & ~n9748;
  assign n9750 = n9749 ^ x737;
  assign n9751 = ~x962 & ~n9750;
  assign n9752 = n8777 ^ x738;
  assign n9753 = n9752 ^ x738;
  assign n9754 = x1121 ^ x738;
  assign n9755 = n9753 & ~n9754;
  assign n9756 = n9755 ^ x738;
  assign n9757 = ~x962 & ~n9756;
  assign n9758 = ~x952 & n7635;
  assign n9759 = n9758 ^ x739;
  assign n9760 = n9759 ^ x739;
  assign n9761 = x1108 ^ x739;
  assign n9762 = n9760 & n9761;
  assign n9763 = n9762 ^ x739;
  assign n9764 = ~x966 & ~n9763;
  assign n9765 = n9758 ^ x741;
  assign n9766 = n9765 ^ x741;
  assign n9767 = x1114 ^ x741;
  assign n9768 = n9766 & ~n9767;
  assign n9769 = n9768 ^ x741;
  assign n9770 = ~x966 & n9769;
  assign n9771 = n9758 ^ x742;
  assign n9772 = n9771 ^ x742;
  assign n9773 = x1112 ^ x742;
  assign n9774 = n9772 & ~n9773;
  assign n9775 = n9774 ^ x742;
  assign n9776 = ~x966 & n9775;
  assign n9777 = n9758 ^ x743;
  assign n9778 = n9777 ^ x743;
  assign n9779 = x1109 ^ x743;
  assign n9780 = n9778 & n9779;
  assign n9781 = n9780 ^ x743;
  assign n9782 = ~x966 & ~n9781;
  assign n9783 = n9758 ^ x744;
  assign n9784 = n9783 ^ x744;
  assign n9785 = x1131 ^ x744;
  assign n9786 = n9784 & ~n9785;
  assign n9787 = n9786 ^ x744;
  assign n9788 = ~x966 & n9787;
  assign n9789 = n9758 ^ x745;
  assign n9790 = n9789 ^ x745;
  assign n9791 = x1111 ^ x745;
  assign n9792 = n9790 & ~n9791;
  assign n9793 = n9792 ^ x745;
  assign n9794 = ~x966 & n9793;
  assign n9795 = n9758 ^ x746;
  assign n9796 = n9795 ^ x746;
  assign n9797 = x1104 ^ x746;
  assign n9798 = n9796 & n9797;
  assign n9799 = n9798 ^ x746;
  assign n9800 = ~x966 & ~n9799;
  assign n9801 = x773 & n9672;
  assign n9802 = n9801 ^ x747;
  assign n9803 = ~n9574 & n9802;
  assign n9804 = n9758 ^ x748;
  assign n9805 = n9804 ^ x748;
  assign n9806 = x1106 ^ x748;
  assign n9807 = n9805 & n9806;
  assign n9808 = n9807 ^ x748;
  assign n9809 = ~x966 & ~n9808;
  assign n9810 = n9758 ^ x749;
  assign n9811 = n9810 ^ x749;
  assign n9812 = x1105 ^ x749;
  assign n9813 = n9811 & n9812;
  assign n9814 = n9813 ^ x749;
  assign n9815 = ~x966 & ~n9814;
  assign n9816 = n9758 ^ x750;
  assign n9817 = n9816 ^ x750;
  assign n9818 = x1130 ^ x750;
  assign n9819 = n9817 & ~n9818;
  assign n9820 = n9819 ^ x750;
  assign n9821 = ~x966 & n9820;
  assign n9822 = n9758 ^ x751;
  assign n9823 = n9822 ^ x751;
  assign n9824 = x1123 ^ x751;
  assign n9825 = n9823 & ~n9824;
  assign n9826 = n9825 ^ x751;
  assign n9827 = ~x966 & n9826;
  assign n9828 = n9758 ^ x752;
  assign n9829 = n9828 ^ x752;
  assign n9830 = x1124 ^ x752;
  assign n9831 = n9829 & ~n9830;
  assign n9832 = n9831 ^ x752;
  assign n9833 = ~x966 & n9832;
  assign n9834 = n9758 ^ x753;
  assign n9835 = n9834 ^ x753;
  assign n9836 = x1117 ^ x753;
  assign n9837 = n9835 & ~n9836;
  assign n9838 = n9837 ^ x753;
  assign n9839 = ~x966 & n9838;
  assign n9840 = n9758 ^ x754;
  assign n9841 = n9840 ^ x754;
  assign n9842 = x1118 ^ x754;
  assign n9843 = n9841 & ~n9842;
  assign n9844 = n9843 ^ x754;
  assign n9845 = ~x966 & n9844;
  assign n9846 = n9758 ^ x755;
  assign n9847 = n9846 ^ x755;
  assign n9848 = x1120 ^ x755;
  assign n9849 = n9847 & ~n9848;
  assign n9850 = n9849 ^ x755;
  assign n9851 = ~x966 & n9850;
  assign n9852 = n9758 ^ x756;
  assign n9853 = n9852 ^ x756;
  assign n9854 = x1119 ^ x756;
  assign n9855 = n9853 & ~n9854;
  assign n9856 = n9855 ^ x756;
  assign n9857 = ~x966 & n9856;
  assign n9858 = n9758 ^ x757;
  assign n9859 = n9858 ^ x757;
  assign n9860 = x1113 ^ x757;
  assign n9861 = n9859 & ~n9860;
  assign n9862 = n9861 ^ x757;
  assign n9863 = ~x966 & n9862;
  assign n9864 = n9758 ^ x758;
  assign n9865 = n9864 ^ x758;
  assign n9866 = x1101 ^ x758;
  assign n9867 = n9865 & n9866;
  assign n9868 = n9867 ^ x758;
  assign n9869 = ~x966 & ~n9868;
  assign n9870 = n9758 ^ x759;
  assign n9871 = n9870 ^ x759;
  assign n9872 = x1100 ^ x759;
  assign n9873 = n9871 & n9872;
  assign n9874 = n9873 ^ x759;
  assign n9875 = ~x966 & ~n9874;
  assign n9876 = n9758 ^ x760;
  assign n9877 = n9876 ^ x760;
  assign n9878 = x1115 ^ x760;
  assign n9879 = n9877 & ~n9878;
  assign n9880 = n9879 ^ x760;
  assign n9881 = ~x966 & n9880;
  assign n9882 = n9758 ^ x761;
  assign n9883 = n9882 ^ x761;
  assign n9884 = x1121 ^ x761;
  assign n9885 = n9883 & ~n9884;
  assign n9886 = n9885 ^ x761;
  assign n9887 = ~x966 & n9886;
  assign n9888 = n9758 ^ x762;
  assign n9889 = n9888 ^ x762;
  assign n9890 = x1129 ^ x762;
  assign n9891 = n9889 & ~n9890;
  assign n9892 = n9891 ^ x762;
  assign n9893 = ~x966 & n9892;
  assign n9894 = n9758 ^ x763;
  assign n9895 = n9894 ^ x763;
  assign n9896 = x1103 ^ x763;
  assign n9897 = n9895 & n9896;
  assign n9898 = n9897 ^ x763;
  assign n9899 = ~x966 & ~n9898;
  assign n9900 = n9758 ^ x764;
  assign n9901 = n9900 ^ x764;
  assign n9902 = x1107 ^ x764;
  assign n9903 = n9901 & n9902;
  assign n9904 = n9903 ^ x764;
  assign n9905 = ~x966 & ~n9904;
  assign n9906 = ~x773 & ~x794;
  assign n9907 = ~x795 & ~x816;
  assign n9908 = n9906 & n9907;
  assign n9909 = ~x721 & ~x747;
  assign n9910 = ~x765 & ~x771;
  assign n9911 = n9909 & n9910;
  assign n9912 = n9908 & n9911;
  assign n9913 = n9574 & ~n9912;
  assign n9914 = x945 ^ x765;
  assign n9915 = ~n9913 & ~n9914;
  assign n9916 = n9758 ^ x766;
  assign n9917 = n9916 ^ x766;
  assign n9918 = x1110 ^ x766;
  assign n9919 = n9917 & n9918;
  assign n9920 = n9919 ^ x766;
  assign n9921 = ~x966 & ~n9920;
  assign n9922 = n9758 ^ x767;
  assign n9923 = n9922 ^ x767;
  assign n9924 = x1116 ^ x767;
  assign n9925 = n9923 & ~n9924;
  assign n9926 = n9925 ^ x767;
  assign n9927 = ~x966 & n9926;
  assign n9928 = n9758 ^ x768;
  assign n9929 = n9928 ^ x768;
  assign n9930 = x1125 ^ x768;
  assign n9931 = n9929 & ~n9930;
  assign n9932 = n9931 ^ x768;
  assign n9933 = ~x966 & n9932;
  assign n9934 = n9557 ^ x769;
  assign n9935 = ~n9574 & n9934;
  assign n9936 = n9758 ^ x770;
  assign n9937 = n9936 ^ x770;
  assign n9938 = x1126 ^ x770;
  assign n9939 = n9937 & ~n9938;
  assign n9940 = n9939 ^ x770;
  assign n9941 = ~x966 & n9940;
  assign n9942 = x987 ^ x771;
  assign n9943 = ~x945 & n9942;
  assign n9944 = n9943 ^ x771;
  assign n9945 = ~n9913 & n9944;
  assign n9946 = n9758 ^ x772;
  assign n9947 = n9946 ^ x772;
  assign n9948 = x1102 ^ x772;
  assign n9949 = n9947 & n9948;
  assign n9950 = n9949 ^ x772;
  assign n9951 = ~x966 & ~n9950;
  assign n9952 = n9672 ^ x773;
  assign n9953 = ~n9913 & n9952;
  assign n9954 = n9758 ^ x774;
  assign n9955 = n9954 ^ x774;
  assign n9956 = x1127 ^ x774;
  assign n9957 = n9955 & ~n9956;
  assign n9958 = n9957 ^ x774;
  assign n9959 = ~x966 & n9958;
  assign n9960 = x765 & x771;
  assign n9961 = n9555 & n9960;
  assign n9962 = n9961 ^ x775;
  assign n9963 = ~n9574 & n9962;
  assign n9964 = n9758 ^ x776;
  assign n9965 = n9964 ^ x776;
  assign n9966 = x1128 ^ x776;
  assign n9967 = n9965 & ~n9966;
  assign n9968 = n9967 ^ x776;
  assign n9969 = ~x966 & n9968;
  assign n9970 = n9758 ^ x777;
  assign n9971 = n9970 ^ x777;
  assign n9972 = x1122 ^ x777;
  assign n9973 = n9971 & ~n9972;
  assign n9974 = n9973 ^ x777;
  assign n9975 = ~x966 & n9974;
  assign n9976 = x832 & x956;
  assign n9977 = ~x1083 & x1085;
  assign n9978 = n9976 & n9977;
  assign n9979 = ~x1046 & n9978;
  assign n9980 = ~x968 & n9979;
  assign n9981 = x1100 ^ x778;
  assign n9982 = n9980 & n9981;
  assign n9983 = n9982 ^ x778;
  assign n9984 = x779 & ~n7717;
  assign n9985 = x780 & ~n7613;
  assign n9986 = x1101 ^ x781;
  assign n9987 = n9980 & n9986;
  assign n9988 = n9987 ^ x781;
  assign n9989 = ~n2380 & ~n7651;
  assign n9990 = ~n7612 & n9989;
  assign n9991 = x1109 ^ x783;
  assign n9992 = n9980 & n9991;
  assign n9993 = n9992 ^ x783;
  assign n9994 = x1110 ^ x784;
  assign n9995 = n9980 & n9994;
  assign n9996 = n9995 ^ x784;
  assign n9997 = x1102 ^ x785;
  assign n9998 = n9980 & n9997;
  assign n9999 = n9998 ^ x785;
  assign n10000 = x786 ^ x24;
  assign n10001 = x954 & n10000;
  assign n10002 = n10001 ^ x24;
  assign n10003 = x1104 ^ x787;
  assign n10004 = n9980 & n10003;
  assign n10005 = n10004 ^ x787;
  assign n10006 = x1105 ^ x788;
  assign n10007 = n9980 & n10006;
  assign n10008 = n10007 ^ x788;
  assign n10009 = x1106 ^ x789;
  assign n10010 = n9980 & n10009;
  assign n10011 = n10010 ^ x789;
  assign n10012 = x1107 ^ x790;
  assign n10013 = n9980 & n10012;
  assign n10014 = n10013 ^ x790;
  assign n10015 = x1108 ^ x791;
  assign n10016 = n9980 & n10015;
  assign n10017 = n10016 ^ x791;
  assign n10018 = x1103 ^ x792;
  assign n10019 = n9980 & n10018;
  assign n10020 = n10019 ^ x792;
  assign n10021 = x968 & n9979;
  assign n10022 = x1130 ^ x794;
  assign n10023 = n10021 & n10022;
  assign n10024 = n10023 ^ x794;
  assign n10025 = x1128 ^ x795;
  assign n10026 = n10021 & n10025;
  assign n10027 = n10026 ^ x795;
  assign n10028 = x266 & ~x269;
  assign n10029 = x279 & n10028;
  assign n10030 = x278 & ~x280;
  assign n10031 = n10029 & n10030;
  assign n10032 = n7996 & n7998;
  assign n10033 = n10031 & n10032;
  assign n10034 = n10033 ^ x264;
  assign n10035 = x1124 ^ x798;
  assign n10036 = n10021 & n10035;
  assign n10037 = n10036 ^ x798;
  assign n10038 = x1107 ^ x799;
  assign n10039 = n10021 & ~n10038;
  assign n10040 = n10039 ^ x799;
  assign n10041 = x1125 ^ x800;
  assign n10042 = n10021 & n10041;
  assign n10043 = n10042 ^ x800;
  assign n10044 = x1126 ^ x801;
  assign n10045 = n10021 & n10044;
  assign n10046 = n10045 ^ x801;
  assign n10047 = ~x274 & n8001;
  assign n10048 = x1106 ^ x803;
  assign n10049 = n10021 & ~n10048;
  assign n10050 = n10049 ^ x803;
  assign n10051 = x1109 ^ x804;
  assign n10052 = n10021 & n10051;
  assign n10053 = n10052 ^ x804;
  assign n10054 = n7997 ^ x270;
  assign n10055 = x1127 ^ x807;
  assign n10056 = n10021 & n10055;
  assign n10057 = n10056 ^ x807;
  assign n10058 = x1101 ^ x808;
  assign n10059 = n10021 & n10058;
  assign n10060 = n10059 ^ x808;
  assign n10061 = x1103 ^ x809;
  assign n10062 = n10021 & ~n10061;
  assign n10063 = n10062 ^ x809;
  assign n10064 = x1108 ^ x810;
  assign n10065 = n10021 & n10064;
  assign n10066 = n10065 ^ x810;
  assign n10067 = x1102 ^ x811;
  assign n10068 = n10021 & n10067;
  assign n10069 = n10068 ^ x811;
  assign n10070 = x1104 ^ x812;
  assign n10071 = n10021 & ~n10070;
  assign n10072 = n10071 ^ x812;
  assign n10073 = x1131 ^ x813;
  assign n10074 = n10021 & n10073;
  assign n10075 = n10074 ^ x813;
  assign n10076 = x1105 ^ x814;
  assign n10077 = n10021 & ~n10076;
  assign n10078 = n10077 ^ x814;
  assign n10079 = x1110 ^ x815;
  assign n10080 = n10021 & n10079;
  assign n10081 = n10080 ^ x815;
  assign n10082 = x1129 ^ x816;
  assign n10083 = n10021 & n10082;
  assign n10084 = n10083 ^ x816;
  assign n10085 = n7994 ^ x269;
  assign n10086 = ~n4056 & ~n4060;
  assign n10087 = n8000 ^ x265;
  assign n10088 = ~x270 & n7997;
  assign n10089 = n10088 ^ x277;
  assign n10090 = ~x811 & ~x893;
  assign n10091 = n1474 & n2872;
  assign n10092 = ~x982 & ~n1473;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = n1476 & ~n10093;
  assign n10095 = x123 & n1537;
  assign n10100 = x1131 ^ x1130;
  assign n10099 = x1129 ^ x1128;
  assign n10101 = n10100 ^ n10099;
  assign n10097 = x1125 ^ x1124;
  assign n10096 = x1127 ^ x1126;
  assign n10098 = n10097 ^ n10096;
  assign n10102 = n10101 ^ n10098;
  assign n10103 = n10102 ^ x825;
  assign n10104 = ~n10095 & ~n10103;
  assign n10105 = n10104 ^ x825;
  assign n10110 = x1123 ^ x1122;
  assign n10109 = x1121 ^ x1120;
  assign n10111 = n10110 ^ n10109;
  assign n10107 = x1117 ^ x1116;
  assign n10106 = x1119 ^ x1118;
  assign n10108 = n10107 ^ n10106;
  assign n10112 = n10111 ^ n10108;
  assign n10113 = n10112 ^ x826;
  assign n10114 = ~n10095 & ~n10113;
  assign n10115 = n10114 ^ x826;
  assign n10120 = x1107 ^ x1106;
  assign n10119 = x1105 ^ x1104;
  assign n10121 = n10120 ^ n10119;
  assign n10117 = x1103 ^ x1102;
  assign n10116 = x1101 ^ x1100;
  assign n10118 = n10117 ^ n10116;
  assign n10122 = n10121 ^ n10118;
  assign n10123 = n10122 ^ x827;
  assign n10124 = ~n10095 & ~n10123;
  assign n10125 = n10124 ^ x827;
  assign n10130 = x1109 ^ x1108;
  assign n10129 = x1111 ^ x1110;
  assign n10131 = n10130 ^ n10129;
  assign n10127 = x1113 ^ x1112;
  assign n10126 = x1115 ^ x1114;
  assign n10128 = n10127 ^ n10126;
  assign n10132 = n10131 ^ n10128;
  assign n10133 = n10132 ^ x828;
  assign n10134 = ~n10095 & ~n10133;
  assign n10135 = n10134 ^ x828;
  assign n10136 = x1091 & n2868;
  assign n10137 = n2872 & n10136;
  assign n10138 = ~x951 & x1092;
  assign n10139 = ~n10137 & ~n10138;
  assign n10140 = n10031 ^ x281;
  assign n10141 = ~x832 & ~x1163;
  assign n10142 = n2907 & n10141;
  assign n10143 = n10136 & n10142;
  assign n10144 = x1091 ^ x833;
  assign n10145 = n2868 & n10144;
  assign n10146 = n10145 ^ x833;
  assign n10147 = x946 & n2868;
  assign n10148 = ~x281 & n7995;
  assign n10149 = n10148 ^ x282;
  assign n10150 = x1049 ^ x837;
  assign n10151 = ~x955 & n10150;
  assign n10152 = n10151 ^ x837;
  assign n10153 = x1047 ^ x838;
  assign n10154 = ~x955 & n10153;
  assign n10155 = n10154 ^ x838;
  assign n10156 = x1074 ^ x839;
  assign n10157 = ~x955 & n10156;
  assign n10158 = n10157 ^ x839;
  assign n10159 = x1196 ^ x840;
  assign n10160 = n2868 & n10159;
  assign n10161 = n10160 ^ x840;
  assign n10162 = x1035 ^ x842;
  assign n10163 = ~x955 & n10162;
  assign n10164 = n10163 ^ x842;
  assign n10165 = x1079 ^ x843;
  assign n10166 = ~x955 & n10165;
  assign n10167 = n10166 ^ x843;
  assign n10168 = x1078 ^ x844;
  assign n10169 = ~x955 & n10168;
  assign n10170 = n10169 ^ x844;
  assign n10171 = x1043 ^ x845;
  assign n10172 = ~x955 & n10171;
  assign n10173 = n10172 ^ x845;
  assign n10174 = x1134 ^ x846;
  assign n10175 = ~n6154 & n10174;
  assign n10176 = n10175 ^ x846;
  assign n10177 = x1055 ^ x847;
  assign n10178 = ~x955 & n10177;
  assign n10179 = n10178 ^ x847;
  assign n10180 = x1039 ^ x848;
  assign n10181 = ~x955 & n10180;
  assign n10182 = n10181 ^ x848;
  assign n10183 = x1198 ^ x849;
  assign n10184 = n2868 & n10183;
  assign n10185 = n10184 ^ x849;
  assign n10186 = x1048 ^ x850;
  assign n10187 = ~x955 & n10186;
  assign n10188 = n10187 ^ x850;
  assign n10189 = x1045 ^ x851;
  assign n10190 = ~x955 & n10189;
  assign n10191 = n10190 ^ x851;
  assign n10192 = x1062 ^ x852;
  assign n10193 = ~x955 & n10192;
  assign n10194 = n10193 ^ x852;
  assign n10195 = x1080 ^ x853;
  assign n10196 = ~x955 & n10195;
  assign n10197 = n10196 ^ x853;
  assign n10198 = x1051 ^ x854;
  assign n10199 = ~x955 & n10198;
  assign n10200 = n10199 ^ x854;
  assign n10201 = x1065 ^ x855;
  assign n10202 = ~x955 & n10201;
  assign n10203 = n10202 ^ x855;
  assign n10204 = x1067 ^ x856;
  assign n10205 = ~x955 & n10204;
  assign n10206 = n10205 ^ x856;
  assign n10207 = x1058 ^ x857;
  assign n10208 = ~x955 & n10207;
  assign n10209 = n10208 ^ x857;
  assign n10210 = x1087 ^ x858;
  assign n10211 = ~x955 & n10210;
  assign n10212 = n10211 ^ x858;
  assign n10213 = x1070 ^ x859;
  assign n10214 = ~x955 & n10213;
  assign n10215 = n10214 ^ x859;
  assign n10216 = x1076 ^ x860;
  assign n10217 = ~x955 & n10216;
  assign n10218 = n10217 ^ x860;
  assign n10219 = x1141 ^ x861;
  assign n10220 = ~n6154 & n10219;
  assign n10221 = n10220 ^ x861;
  assign n10222 = x1139 ^ x862;
  assign n10223 = ~n6154 & n10222;
  assign n10224 = n10223 ^ x862;
  assign n10225 = x1199 ^ x863;
  assign n10226 = n2868 & n10225;
  assign n10227 = n10226 ^ x863;
  assign n10228 = x1197 ^ x864;
  assign n10229 = n2868 & n10228;
  assign n10230 = n10229 ^ x864;
  assign n10231 = x1040 ^ x865;
  assign n10232 = ~x955 & n10231;
  assign n10233 = n10232 ^ x865;
  assign n10234 = x1053 ^ x866;
  assign n10235 = ~x955 & n10234;
  assign n10236 = n10235 ^ x866;
  assign n10237 = x1057 ^ x867;
  assign n10238 = ~x955 & n10237;
  assign n10239 = n10238 ^ x867;
  assign n10240 = x1063 ^ x868;
  assign n10241 = ~x955 & n10240;
  assign n10242 = n10241 ^ x868;
  assign n10243 = x1140 ^ x869;
  assign n10244 = ~n6154 & n10243;
  assign n10245 = n10244 ^ x869;
  assign n10246 = x1069 ^ x870;
  assign n10247 = ~x955 & n10246;
  assign n10248 = n10247 ^ x870;
  assign n10249 = x1072 ^ x871;
  assign n10250 = ~x955 & n10249;
  assign n10251 = n10250 ^ x871;
  assign n10252 = x1084 ^ x872;
  assign n10253 = ~x955 & n10252;
  assign n10254 = n10253 ^ x872;
  assign n10255 = x1044 ^ x873;
  assign n10256 = ~x955 & n10255;
  assign n10257 = n10256 ^ x873;
  assign n10258 = x1036 ^ x874;
  assign n10259 = ~x955 & n10258;
  assign n10260 = n10259 ^ x874;
  assign n10261 = x1136 ^ x875;
  assign n10262 = ~n6154 & n10261;
  assign n10263 = n10262 ^ x875;
  assign n10264 = x1037 ^ x876;
  assign n10265 = ~x955 & n10264;
  assign n10266 = n10265 ^ x876;
  assign n10267 = x1138 ^ x877;
  assign n10268 = ~n6154 & n10267;
  assign n10269 = n10268 ^ x877;
  assign n10270 = x1137 ^ x878;
  assign n10271 = ~n6154 & n10270;
  assign n10272 = n10271 ^ x878;
  assign n10273 = x1135 ^ x879;
  assign n10274 = ~n6154 & n10273;
  assign n10275 = n10274 ^ x879;
  assign n10276 = x1081 ^ x880;
  assign n10277 = ~x955 & n10276;
  assign n10278 = n10277 ^ x880;
  assign n10279 = x1059 ^ x881;
  assign n10280 = ~x955 & n10279;
  assign n10281 = n10280 ^ x881;
  assign n10282 = x1107 ^ x883;
  assign n10283 = ~n10095 & ~n10282;
  assign n10284 = n10283 ^ x883;
  assign n10285 = x1124 ^ x884;
  assign n10286 = ~n10095 & ~n10285;
  assign n10287 = n10286 ^ x884;
  assign n10288 = x1125 ^ x885;
  assign n10289 = ~n10095 & ~n10288;
  assign n10290 = n10289 ^ x885;
  assign n10291 = x1109 ^ x886;
  assign n10292 = ~n10095 & ~n10291;
  assign n10293 = n10292 ^ x886;
  assign n10294 = x1100 ^ x887;
  assign n10295 = ~n10095 & ~n10294;
  assign n10296 = n10295 ^ x887;
  assign n10297 = x1120 ^ x888;
  assign n10298 = ~n10095 & ~n10297;
  assign n10299 = n10298 ^ x888;
  assign n10300 = x1103 ^ x889;
  assign n10301 = ~n10095 & ~n10300;
  assign n10302 = n10301 ^ x889;
  assign n10303 = x1126 ^ x890;
  assign n10304 = ~n10095 & ~n10303;
  assign n10305 = n10304 ^ x890;
  assign n10306 = x1116 ^ x891;
  assign n10307 = ~n10095 & ~n10306;
  assign n10308 = n10307 ^ x891;
  assign n10309 = x1101 ^ x892;
  assign n10310 = ~n10095 & ~n10309;
  assign n10311 = n10310 ^ x892;
  assign n10312 = x1119 ^ x894;
  assign n10313 = ~n10095 & ~n10312;
  assign n10314 = n10313 ^ x894;
  assign n10315 = x1113 ^ x895;
  assign n10316 = ~n10095 & ~n10315;
  assign n10317 = n10316 ^ x895;
  assign n10318 = x1118 ^ x896;
  assign n10319 = ~n10095 & ~n10318;
  assign n10320 = n10319 ^ x896;
  assign n10321 = x1129 ^ x898;
  assign n10322 = ~n10095 & ~n10321;
  assign n10323 = n10322 ^ x898;
  assign n10324 = x1115 ^ x899;
  assign n10325 = ~n10095 & ~n10324;
  assign n10326 = n10325 ^ x899;
  assign n10327 = x1110 ^ x900;
  assign n10328 = ~n10095 & ~n10327;
  assign n10329 = n10328 ^ x900;
  assign n10330 = x1111 ^ x902;
  assign n10331 = ~n10095 & ~n10330;
  assign n10332 = n10331 ^ x902;
  assign n10333 = x1121 ^ x903;
  assign n10334 = ~n10095 & ~n10333;
  assign n10335 = n10334 ^ x903;
  assign n10336 = x1127 ^ x904;
  assign n10337 = ~n10095 & ~n10336;
  assign n10338 = n10337 ^ x904;
  assign n10339 = x1131 ^ x905;
  assign n10340 = ~n10095 & ~n10339;
  assign n10341 = n10340 ^ x905;
  assign n10342 = x1128 ^ x906;
  assign n10343 = ~n10095 & ~n10342;
  assign n10344 = n10343 ^ x906;
  assign n10345 = ~x624 & ~x979;
  assign n10346 = x604 & n10345;
  assign n10347 = ~x598 & x979;
  assign n10348 = ~x615 & n10347;
  assign n10349 = ~n10346 & ~n10348;
  assign n10350 = n10349 ^ x907;
  assign n10351 = x782 & ~n10350;
  assign n10352 = n10351 ^ x907;
  assign n10353 = x1122 ^ x908;
  assign n10354 = ~n10095 & ~n10353;
  assign n10355 = n10354 ^ x908;
  assign n10356 = x1105 ^ x909;
  assign n10357 = ~n10095 & ~n10356;
  assign n10358 = n10357 ^ x909;
  assign n10359 = x1117 ^ x910;
  assign n10360 = ~n10095 & ~n10359;
  assign n10361 = n10360 ^ x910;
  assign n10362 = x1130 ^ x911;
  assign n10363 = ~n10095 & ~n10362;
  assign n10364 = n10363 ^ x911;
  assign n10365 = x1114 ^ x912;
  assign n10366 = ~n10095 & ~n10365;
  assign n10367 = n10366 ^ x912;
  assign n10368 = x1106 ^ x913;
  assign n10369 = ~n10095 & ~n10368;
  assign n10370 = n10369 ^ x913;
  assign n10371 = n7993 ^ x280;
  assign n10372 = x1108 ^ x915;
  assign n10373 = ~n10095 & ~n10372;
  assign n10374 = n10373 ^ x915;
  assign n10375 = x1123 ^ x916;
  assign n10376 = ~n10095 & ~n10375;
  assign n10377 = n10376 ^ x916;
  assign n10378 = x1112 ^ x917;
  assign n10379 = ~n10095 & ~n10378;
  assign n10380 = n10379 ^ x917;
  assign n10381 = x1104 ^ x918;
  assign n10382 = ~n10095 & ~n10381;
  assign n10383 = n10382 ^ x918;
  assign n10384 = x1102 ^ x919;
  assign n10385 = ~n10095 & ~n10384;
  assign n10386 = n10385 ^ x919;
  assign n10387 = x1139 ^ x920;
  assign n10388 = x1093 & n10387;
  assign n10389 = n10388 ^ x920;
  assign n10390 = x1140 ^ x921;
  assign n10391 = x1093 & n10390;
  assign n10392 = n10391 ^ x921;
  assign n10393 = x1152 ^ x922;
  assign n10394 = x1093 & n10393;
  assign n10395 = n10394 ^ x922;
  assign n10396 = x1154 ^ x923;
  assign n10397 = x1093 & n10396;
  assign n10398 = n10397 ^ x923;
  assign n10399 = x311 & n6507;
  assign n10400 = x1155 ^ x925;
  assign n10401 = x1093 & n10400;
  assign n10402 = n10401 ^ x925;
  assign n10403 = x1157 ^ x926;
  assign n10404 = x1093 & n10403;
  assign n10405 = n10404 ^ x926;
  assign n10406 = x1145 ^ x927;
  assign n10407 = x1093 & n10406;
  assign n10408 = n10407 ^ x927;
  assign n10409 = x1136 ^ x928;
  assign n10410 = x1093 & n10409;
  assign n10411 = n10410 ^ x928;
  assign n10412 = x1144 ^ x929;
  assign n10413 = x1093 & n10412;
  assign n10414 = n10413 ^ x929;
  assign n10415 = x1134 ^ x930;
  assign n10416 = x1093 & n10415;
  assign n10417 = n10416 ^ x930;
  assign n10418 = x1150 ^ x931;
  assign n10419 = x1093 & n10418;
  assign n10420 = n10419 ^ x931;
  assign n10421 = x1093 & n1855;
  assign n10422 = n10421 ^ x932;
  assign n10423 = x1137 ^ x933;
  assign n10424 = x1093 & n10423;
  assign n10425 = n10424 ^ x933;
  assign n10426 = x1147 ^ x934;
  assign n10427 = x1093 & n10426;
  assign n10428 = n10427 ^ x934;
  assign n10429 = x1141 ^ x935;
  assign n10430 = x1093 & n10429;
  assign n10431 = n10430 ^ x935;
  assign n10432 = x1149 ^ x936;
  assign n10433 = x1093 & n10432;
  assign n10434 = n10433 ^ x936;
  assign n10435 = x1148 ^ x937;
  assign n10436 = x1093 & n10435;
  assign n10437 = n10436 ^ x937;
  assign n10438 = x1135 ^ x938;
  assign n10439 = x1093 & n10438;
  assign n10440 = n10439 ^ x938;
  assign n10441 = x1146 ^ x939;
  assign n10442 = x1093 & n10441;
  assign n10443 = n10442 ^ x939;
  assign n10444 = x1138 ^ x940;
  assign n10445 = x1093 & n10444;
  assign n10446 = n10445 ^ x940;
  assign n10447 = x1153 ^ x941;
  assign n10448 = x1093 & n10447;
  assign n10449 = n10448 ^ x941;
  assign n10450 = x1156 ^ x942;
  assign n10451 = x1093 & n10450;
  assign n10452 = n10451 ^ x942;
  assign n10453 = x1151 ^ x943;
  assign n10454 = x1093 & n10453;
  assign n10455 = n10454 ^ x943;
  assign n10456 = x1143 ^ x944;
  assign n10457 = x1093 & n10456;
  assign n10458 = n10457 ^ x944;
  assign n10459 = x230 & n2868;
  assign n10460 = ~n10345 & ~n10347;
  assign n10461 = n10460 ^ x947;
  assign n10462 = x782 & n10461;
  assign n10463 = n10462 ^ x947;
  assign n10464 = x992 ^ x266;
  assign n10465 = x949 ^ x313;
  assign n10466 = x954 & ~n10465;
  assign n10467 = n10466 ^ x313;
  assign n10468 = x1092 & n1473;
  assign n10469 = x957 & x1092;
  assign n10470 = ~x31 & ~n10469;
  assign n10471 = ~x782 & x960;
  assign n10472 = ~x230 & x961;
  assign n10473 = ~x782 & x963;
  assign n10474 = ~x230 & x967;
  assign n10475 = ~x230 & x969;
  assign n10476 = ~x782 & x970;
  assign n10477 = ~x230 & x971;
  assign n10478 = ~x782 & x972;
  assign n10479 = ~x230 & x974;
  assign n10480 = ~x782 & x975;
  assign n10481 = ~x230 & x977;
  assign n10482 = ~x782 & x978;
  assign n10483 = ~x598 & x615;
  assign n10484 = x824 & x1092;
  assign n10485 = ~x604 & ~x624;
  assign y0 = x668;
  assign y1 = x672;
  assign y2 = x664;
  assign y3 = x667;
  assign y4 = x676;
  assign y5 = x673;
  assign y6 = x675;
  assign y7 = x666;
  assign y8 = x679;
  assign y9 = x674;
  assign y10 = x663;
  assign y11 = x670;
  assign y12 = x677;
  assign y13 = x682;
  assign y14 = x671;
  assign y15 = x678;
  assign y16 = x718;
  assign y17 = x707;
  assign y18 = x708;
  assign y19 = x713;
  assign y20 = x711;
  assign y21 = x716;
  assign y22 = x733;
  assign y23 = x712;
  assign y24 = x689;
  assign y25 = x717;
  assign y26 = x692;
  assign y27 = x719;
  assign y28 = x722;
  assign y29 = x714;
  assign y30 = x720;
  assign y31 = x685;
  assign y32 = x837;
  assign y33 = x850;
  assign y34 = x872;
  assign y35 = x871;
  assign y36 = x881;
  assign y37 = x866;
  assign y38 = x876;
  assign y39 = x873;
  assign y40 = x874;
  assign y41 = x859;
  assign y42 = x855;
  assign y43 = x852;
  assign y44 = x870;
  assign y45 = x848;
  assign y46 = x865;
  assign y47 = x856;
  assign y48 = x853;
  assign y49 = x847;
  assign y50 = x857;
  assign y51 = x854;
  assign y52 = x858;
  assign y53 = x845;
  assign y54 = x838;
  assign y55 = x842;
  assign y56 = x843;
  assign y57 = x839;
  assign y58 = x844;
  assign y59 = x868;
  assign y60 = x851;
  assign y61 = x867;
  assign y62 = x880;
  assign y63 = x860;
  assign y64 = x1030;
  assign y65 = x1034;
  assign y66 = x1015;
  assign y67 = x1020;
  assign y68 = x1025;
  assign y69 = x1005;
  assign y70 = x996;
  assign y71 = x1012;
  assign y72 = x993;
  assign y73 = x1016;
  assign y74 = x1021;
  assign y75 = x1010;
  assign y76 = x1027;
  assign y77 = x1018;
  assign y78 = x1017;
  assign y79 = x1024;
  assign y80 = x1009;
  assign y81 = x1032;
  assign y82 = x1003;
  assign y83 = x997;
  assign y84 = x1013;
  assign y85 = x1011;
  assign y86 = x1008;
  assign y87 = x1019;
  assign y88 = x1031;
  assign y89 = x1022;
  assign y90 = x1000;
  assign y91 = x1023;
  assign y92 = x1002;
  assign y93 = x1026;
  assign y94 = x1006;
  assign y95 = x998;
  assign y96 = x31;
  assign y97 = x80;
  assign y98 = x893;
  assign y99 = x467;
  assign y100 = x78;
  assign y101 = x112;
  assign y102 = x13;
  assign y103 = x25;
  assign y104 = x226;
  assign y105 = x127;
  assign y106 = x822;
  assign y107 = x808;
  assign y108 = x227;
  assign y109 = x477;
  assign y110 = x834;
  assign y111 = x229;
  assign y112 = x12;
  assign y113 = x11;
  assign y114 = x10;
  assign y115 = x9;
  assign y116 = x8;
  assign y117 = x7;
  assign y118 = x6;
  assign y119 = x5;
  assign y120 = x4;
  assign y121 = x3;
  assign y122 = x0;
  assign y123 = x2;
  assign y124 = x1;
  assign y125 = x310;
  assign y126 = x302;
  assign y127 = x475;
  assign y128 = x474;
  assign y129 = x466;
  assign y130 = x473;
  assign y131 = x471;
  assign y132 = x472;
  assign y133 = x470;
  assign y134 = x469;
  assign y135 = x465;
  assign y136 = x1028;
  assign y137 = x1033;
  assign y138 = x995;
  assign y139 = x994;
  assign y140 = x28;
  assign y141 = x27;
  assign y142 = x26;
  assign y143 = x29;
  assign y144 = x15;
  assign y145 = x14;
  assign y146 = x21;
  assign y147 = x20;
  assign y148 = x19;
  assign y149 = x18;
  assign y150 = x17;
  assign y151 = x16;
  assign y152 = x1096;
  assign y153 = ~n1734;
  assign y154 = ~n1785;
  assign y155 = ~n1805;
  assign y156 = ~n1850;
  assign y157 = ~n1919;
  assign y158 = n1966;
  assign y159 = ~n2024;
  assign y160 = ~n2070;
  assign y161 = n2115;
  assign y162 = n2175;
  assign y163 = n2222;
  assign y164 = n2259;
  assign y165 = n2296;
  assign y166 = ~1'b0;
  assign y167 = ~n2411;
  assign y168 = x228;
  assign y169 = x22;
  assign y170 = ~x1090;
  assign y171 = n2514;
  assign y172 = n2522;
  assign y173 = n2526;
  assign y174 = ~n2540;
  assign y175 = n2543;
  assign y176 = n2546;
  assign y177 = n2549;
  assign y178 = n2552;
  assign y179 = x1089;
  assign y180 = x23;
  assign y181 = ~n2411;
  assign y182 = ~n2580;
  assign y183 = n2586;
  assign y184 = n2592;
  assign y185 = n2594;
  assign y186 = n2596;
  assign y187 = n2598;
  assign y188 = x37;
  assign y189 = ~n2911;
  assign y190 = ~n2944;
  assign y191 = ~n3104;
  assign y192 = n3204;
  assign y193 = n3257;
  assign y194 = n3263;
  assign y195 = ~n2577;
  assign y196 = ~n3275;
  assign y197 = ~n3309;
  assign y198 = n3314;
  assign y199 = n3364;
  assign y200 = ~n3397;
  assign y201 = ~n3412;
  assign y202 = ~n3419;
  assign y203 = n3420;
  assign y204 = ~n3427;
  assign y205 = n3441;
  assign y206 = n3443;
  assign y207 = ~n3447;
  assign y208 = ~n3466;
  assign y209 = n3471;
  assign y210 = ~n3489;
  assign y211 = ~n3497;
  assign y212 = ~n3501;
  assign y213 = ~n3504;
  assign y214 = n3511;
  assign y215 = ~n3516;
  assign y216 = n3518;
  assign y217 = ~n3523;
  assign y218 = ~n3529;
  assign y219 = ~n3532;
  assign y220 = n3537;
  assign y221 = ~n3541;
  assign y222 = ~n3544;
  assign y223 = n3546;
  assign y224 = n3555;
  assign y225 = n3560;
  assign y226 = n3566;
  assign y227 = n3569;
  assign y228 = ~n3584;
  assign y229 = ~n3595;
  assign y230 = ~n3604;
  assign y231 = n3610;
  assign y232 = ~n3621;
  assign y233 = ~n3624;
  assign y234 = n3637;
  assign y235 = n3640;
  assign y236 = n3641;
  assign y237 = ~n3749;
  assign y238 = n3778;
  assign y239 = n3781;
  assign y240 = n3785;
  assign y241 = ~n3791;
  assign y242 = n3795;
  assign y243 = n3798;
  assign y244 = n3799;
  assign y245 = n3800;
  assign y246 = ~n3806;
  assign y247 = n3810;
  assign y248 = ~n3813;
  assign y249 = ~n3824;
  assign y250 = n3833;
  assign y251 = ~n3837;
  assign y252 = ~n3841;
  assign y253 = ~n3853;
  assign y254 = n3868;
  assign y255 = ~n3873;
  assign y256 = n3876;
  assign y257 = ~n3886;
  assign y258 = n3896;
  assign y259 = ~n3903;
  assign y260 = n3904;
  assign y261 = n3905;
  assign y262 = ~n3910;
  assign y263 = x117;
  assign y264 = ~n3913;
  assign y265 = n3914;
  assign y266 = ~n3919;
  assign y267 = n3920;
  assign y268 = ~n3924;
  assign y269 = ~n3928;
  assign y270 = ~n3929;
  assign y271 = n3932;
  assign y272 = n3934;
  assign y273 = n3937;
  assign y274 = n3939;
  assign y275 = ~n2583;
  assign y276 = n4037;
  assign y277 = n4051;
  assign y278 = n4063;
  assign y279 = n4119;
  assign y280 = ~n4054;
  assign y281 = n4132;
  assign y282 = ~n4214;
  assign y283 = n4275;
  assign y284 = n4284;
  assign y285 = x131;
  assign y286 = ~n4293;
  assign y287 = ~n4333;
  assign y288 = ~n4048;
  assign y289 = n4389;
  assign y290 = n4412;
  assign y291 = n4437;
  assign y292 = n4454;
  assign y293 = n4482;
  assign y294 = ~n4489;
  assign y295 = ~n4519;
  assign y296 = ~n4529;
  assign y297 = ~n4617;
  assign y298 = ~n4628;
  assign y299 = n4639;
  assign y300 = ~n4650;
  assign y301 = n4661;
  assign y302 = ~n4672;
  assign y303 = n4681;
  assign y304 = ~n4692;
  assign y305 = ~n4701;
  assign y306 = ~n4721;
  assign y307 = ~n4732;
  assign y308 = ~n4743;
  assign y309 = n4754;
  assign y310 = ~n4765;
  assign y311 = ~n4776;
  assign y312 = ~n4787;
  assign y313 = ~n4798;
  assign y314 = ~n4809;
  assign y315 = ~n4820;
  assign y316 = ~n4831;
  assign y317 = ~n4842;
  assign y318 = n4851;
  assign y319 = ~n4860;
  assign y320 = ~n4871;
  assign y321 = ~n4882;
  assign y322 = ~n4891;
  assign y323 = n4902;
  assign y324 = ~n4913;
  assign y325 = ~n4924;
  assign y326 = ~n4935;
  assign y327 = ~n4946;
  assign y328 = ~n4957;
  assign y329 = ~n4968;
  assign y330 = ~n4977;
  assign y331 = n4986;
  assign y332 = ~n4995;
  assign y333 = ~n5004;
  assign y334 = ~n5013;
  assign y335 = ~n5022;
  assign y336 = ~n5031;
  assign y337 = ~n5040;
  assign y338 = ~n5049;
  assign y339 = ~n5058;
  assign y340 = ~n5067;
  assign y341 = ~n5076;
  assign y342 = ~n5085;
  assign y343 = ~n5094;
  assign y344 = ~n5103;
  assign y345 = ~n5112;
  assign y346 = n5121;
  assign y347 = ~n5130;
  assign y348 = ~n5139;
  assign y349 = ~n5148;
  assign y350 = ~n5157;
  assign y351 = ~n5166;
  assign y352 = ~n5180;
  assign y353 = ~n5194;
  assign y354 = ~n5203;
  assign y355 = n5214;
  assign y356 = n5225;
  assign y357 = n5236;
  assign y358 = ~n5275;
  assign y359 = ~n5283;
  assign y360 = ~n5290;
  assign y361 = ~n5304;
  assign y362 = ~n5308;
  assign y363 = ~n5315;
  assign y364 = ~n5326;
  assign y365 = ~n5337;
  assign y366 = ~n5348;
  assign y367 = n5357;
  assign y368 = n5366;
  assign y369 = ~n5375;
  assign y370 = ~n5384;
  assign y371 = ~n5393;
  assign y372 = n5404;
  assign y373 = n5415;
  assign y374 = ~n5426;
  assign y375 = ~n5430;
  assign y376 = ~n5439;
  assign y377 = ~n5443;
  assign y378 = n5454;
  assign y379 = n5463;
  assign y380 = n5472;
  assign y381 = n5481;
  assign y382 = ~n5491;
  assign y383 = n5500;
  assign y384 = ~n5510;
  assign y385 = ~n5518;
  assign y386 = x232;
  assign y387 = n5522;
  assign y388 = x236;
  assign y389 = ~n5530;
  assign y390 = ~n5660;
  assign y391 = n5700;
  assign y392 = n5739;
  assign y393 = ~n5497;
  assign y394 = n5839;
  assign y395 = n5878;
  assign y396 = n5898;
  assign y397 = n5920;
  assign y398 = n5934;
  assign y399 = n5961;
  assign y400 = ~n5998;
  assign y401 = n6017;
  assign y402 = n6031;
  assign y403 = n6045;
  assign y404 = n6051;
  assign y405 = n6065;
  assign y406 = n6071;
  assign y407 = n6073;
  assign y408 = n6085;
  assign y409 = ~n6091;
  assign y410 = n6100;
  assign y411 = n6109;
  assign y412 = n6115;
  assign y413 = n6121;
  assign y414 = n6127;
  assign y415 = n6133;
  assign y416 = n6139;
  assign y417 = n6145;
  assign y418 = n6151;
  assign y419 = ~n6162;
  assign y420 = ~n6171;
  assign y421 = ~n6182;
  assign y422 = ~n6193;
  assign y423 = n6204;
  assign y424 = n6213;
  assign y425 = n6222;
  assign y426 = ~n6233;
  assign y427 = ~n6244;
  assign y428 = n6253;
  assign y429 = n6262;
  assign y430 = n6271;
  assign y431 = ~n6282;
  assign y432 = n6291;
  assign y433 = n6300;
  assign y434 = ~n6311;
  assign y435 = n6322;
  assign y436 = n6333;
  assign y437 = ~n6344;
  assign y438 = ~n6355;
  assign y439 = ~n6366;
  assign y440 = n6375;
  assign y441 = ~n6384;
  assign y442 = n6396;
  assign y443 = ~n6405;
  assign y444 = n6407;
  assign y445 = n6410;
  assign y446 = n6422;
  assign y447 = n6425;
  assign y448 = n6428;
  assign y449 = n6431;
  assign y450 = n6434;
  assign y451 = n6437;
  assign y452 = n6440;
  assign y453 = n6443;
  assign y454 = n6446;
  assign y455 = n6449;
  assign y456 = ~n6456;
  assign y457 = ~n6460;
  assign y458 = n6464;
  assign y459 = ~n6478;
  assign y460 = n6481;
  assign y461 = n6484;
  assign y462 = n6487;
  assign y463 = n6490;
  assign y464 = n6493;
  assign y465 = n6496;
  assign y466 = n6499;
  assign y467 = ~n6506;
  assign y468 = n6510;
  assign y469 = n6512;
  assign y470 = ~n6523;
  assign y471 = n6525;
  assign y472 = n6529;
  assign y473 = n6532;
  assign y474 = n6536;
  assign y475 = n6540;
  assign y476 = n6543;
  assign y477 = n6546;
  assign y478 = n6549;
  assign y479 = n6552;
  assign y480 = n6555;
  assign y481 = n6558;
  assign y482 = n6561;
  assign y483 = n6564;
  assign y484 = n6567;
  assign y485 = n6570;
  assign y486 = n6573;
  assign y487 = n6578;
  assign y488 = n6582;
  assign y489 = ~n6586;
  assign y490 = n6589;
  assign y491 = n6592;
  assign y492 = n6595;
  assign y493 = n6598;
  assign y494 = n6601;
  assign y495 = n6604;
  assign y496 = n6607;
  assign y497 = ~n6613;
  assign y498 = n6617;
  assign y499 = n6620;
  assign y500 = n6623;
  assign y501 = n6626;
  assign y502 = n6629;
  assign y503 = n6632;
  assign y504 = n6635;
  assign y505 = n6638;
  assign y506 = n6641;
  assign y507 = n6644;
  assign y508 = n6647;
  assign y509 = n6650;
  assign y510 = n6653;
  assign y511 = n6656;
  assign y512 = n6659;
  assign y513 = n6662;
  assign y514 = n6665;
  assign y515 = n6668;
  assign y516 = n6671;
  assign y517 = n6674;
  assign y518 = n6677;
  assign y519 = n6680;
  assign y520 = n6683;
  assign y521 = n6686;
  assign y522 = n6689;
  assign y523 = n6692;
  assign y524 = n6695;
  assign y525 = n6698;
  assign y526 = n6701;
  assign y527 = n6704;
  assign y528 = n6707;
  assign y529 = n6710;
  assign y530 = n6713;
  assign y531 = n6716;
  assign y532 = n6719;
  assign y533 = n6722;
  assign y534 = n6725;
  assign y535 = n6728;
  assign y536 = n6731;
  assign y537 = n6734;
  assign y538 = n6737;
  assign y539 = n6740;
  assign y540 = n6743;
  assign y541 = n6746;
  assign y542 = n6749;
  assign y543 = n6752;
  assign y544 = n6755;
  assign y545 = n6758;
  assign y546 = n6761;
  assign y547 = n6764;
  assign y548 = n6767;
  assign y549 = n6770;
  assign y550 = n6773;
  assign y551 = n6776;
  assign y552 = n6779;
  assign y553 = n6782;
  assign y554 = n6785;
  assign y555 = n6788;
  assign y556 = n6791;
  assign y557 = n6794;
  assign y558 = n6797;
  assign y559 = n6800;
  assign y560 = n6803;
  assign y561 = n6806;
  assign y562 = n6809;
  assign y563 = n6812;
  assign y564 = n6815;
  assign y565 = n6818;
  assign y566 = n6821;
  assign y567 = n6824;
  assign y568 = n6827;
  assign y569 = n6830;
  assign y570 = n6833;
  assign y571 = n6837;
  assign y572 = n6840;
  assign y573 = n6843;
  assign y574 = n6846;
  assign y575 = n6849;
  assign y576 = n6852;
  assign y577 = n6855;
  assign y578 = n6858;
  assign y579 = n6861;
  assign y580 = n6864;
  assign y581 = n6867;
  assign y582 = n6870;
  assign y583 = n6873;
  assign y584 = n6876;
  assign y585 = n6879;
  assign y586 = n6882;
  assign y587 = n6885;
  assign y588 = n6888;
  assign y589 = n6891;
  assign y590 = n6894;
  assign y591 = n6897;
  assign y592 = n6900;
  assign y593 = n6903;
  assign y594 = n6906;
  assign y595 = n6909;
  assign y596 = n6912;
  assign y597 = n6915;
  assign y598 = n6918;
  assign y599 = n6921;
  assign y600 = n6924;
  assign y601 = n6927;
  assign y602 = n6930;
  assign y603 = n6933;
  assign y604 = n6936;
  assign y605 = n6939;
  assign y606 = n6942;
  assign y607 = n6945;
  assign y608 = n6948;
  assign y609 = n6951;
  assign y610 = n6954;
  assign y611 = n6957;
  assign y612 = n6960;
  assign y613 = n6963;
  assign y614 = n6986;
  assign y615 = n6989;
  assign y616 = n6992;
  assign y617 = n6995;
  assign y618 = n6998;
  assign y619 = n7001;
  assign y620 = n7004;
  assign y621 = n7007;
  assign y622 = ~n7012;
  assign y623 = ~n7017;
  assign y624 = ~n7022;
  assign y625 = ~n7025;
  assign y626 = ~n7030;
  assign y627 = ~n7035;
  assign y628 = ~n7040;
  assign y629 = ~n7045;
  assign y630 = ~n7050;
  assign y631 = ~n7055;
  assign y632 = ~n7060;
  assign y633 = ~n7062;
  assign y634 = ~n6520;
  assign y635 = n7063;
  assign y636 = x583;
  assign y637 = n6385;
  assign y638 = n7066;
  assign y639 = n7069;
  assign y640 = n7072;
  assign y641 = n7075;
  assign y642 = n7078;
  assign y643 = n7081;
  assign y644 = n7084;
  assign y645 = n7087;
  assign y646 = n7090;
  assign y647 = n7093;
  assign y648 = n7096;
  assign y649 = n7099;
  assign y650 = n7102;
  assign y651 = n7105;
  assign y652 = n7108;
  assign y653 = n7111;
  assign y654 = n7114;
  assign y655 = n7117;
  assign y656 = n7120;
  assign y657 = n7123;
  assign y658 = n7126;
  assign y659 = n7129;
  assign y660 = n7132;
  assign y661 = n7135;
  assign y662 = n7138;
  assign y663 = n7141;
  assign y664 = n7144;
  assign y665 = n7147;
  assign y666 = n7150;
  assign y667 = n7153;
  assign y668 = n7156;
  assign y669 = n7159;
  assign y670 = n7162;
  assign y671 = n7165;
  assign y672 = n7168;
  assign y673 = n7171;
  assign y674 = n7174;
  assign y675 = n7177;
  assign y676 = n7180;
  assign y677 = n7183;
  assign y678 = n7186;
  assign y679 = n7189;
  assign y680 = n7192;
  assign y681 = n7195;
  assign y682 = n7198;
  assign y683 = n7201;
  assign y684 = n7204;
  assign y685 = n7207;
  assign y686 = n7210;
  assign y687 = n7213;
  assign y688 = n7216;
  assign y689 = n7219;
  assign y690 = n7222;
  assign y691 = n7225;
  assign y692 = n7228;
  assign y693 = n7231;
  assign y694 = n7234;
  assign y695 = n7237;
  assign y696 = n7240;
  assign y697 = n7243;
  assign y698 = n7246;
  assign y699 = n7249;
  assign y700 = n7252;
  assign y701 = n7255;
  assign y702 = n7258;
  assign y703 = n7261;
  assign y704 = n7264;
  assign y705 = n7267;
  assign y706 = n7270;
  assign y707 = n7273;
  assign y708 = n7276;
  assign y709 = n7279;
  assign y710 = n7282;
  assign y711 = n7285;
  assign y712 = n7288;
  assign y713 = n7291;
  assign y714 = n7294;
  assign y715 = n7297;
  assign y716 = n7300;
  assign y717 = n7303;
  assign y718 = n7306;
  assign y719 = n7309;
  assign y720 = n7312;
  assign y721 = n7315;
  assign y722 = n7318;
  assign y723 = n7321;
  assign y724 = n7334;
  assign y725 = n7337;
  assign y726 = n7340;
  assign y727 = n7343;
  assign y728 = n7346;
  assign y729 = n7349;
  assign y730 = n7352;
  assign y731 = n7355;
  assign y732 = n7358;
  assign y733 = n7361;
  assign y734 = n7364;
  assign y735 = n7367;
  assign y736 = n7370;
  assign y737 = n7373;
  assign y738 = n7376;
  assign y739 = n7379;
  assign y740 = ~n2320;
  assign y741 = n7382;
  assign y742 = n7385;
  assign y743 = n7388;
  assign y744 = n7391;
  assign y745 = n7399;
  assign y746 = ~n7424;
  assign y747 = ~n7430;
  assign y748 = n7436;
  assign y749 = n7440;
  assign y750 = ~n7596;
  assign y751 = n7600;
  assign y752 = n7604;
  assign y753 = n7609;
  assign y754 = n7611;
  assign y755 = ~n7617;
  assign y756 = n7620;
  assign y757 = n7622;
  assign y758 = n7628;
  assign y759 = n7631;
  assign y760 = n7649;
  assign y761 = ~n7656;
  assign y762 = n7658;
  assign y763 = n7668;
  assign y764 = n7674;
  assign y765 = n7680;
  assign y766 = n7686;
  assign y767 = n7692;
  assign y768 = n7698;
  assign y769 = n7704;
  assign y770 = n7710;
  assign y771 = n7716;
  assign y772 = ~n7721;
  assign y773 = n7731;
  assign y774 = n7741;
  assign y775 = n7747;
  assign y776 = n7753;
  assign y777 = n7759;
  assign y778 = n7765;
  assign y779 = n7771;
  assign y780 = n7777;
  assign y781 = ~n7783;
  assign y782 = n7794;
  assign y783 = n7800;
  assign y784 = n7806;
  assign y785 = n7812;
  assign y786 = n7818;
  assign y787 = n7824;
  assign y788 = n7830;
  assign y789 = n7836;
  assign y790 = n7842;
  assign y791 = n7848;
  assign y792 = n7854;
  assign y793 = n7860;
  assign y794 = n7866;
  assign y795 = n7872;
  assign y796 = n7878;
  assign y797 = n7884;
  assign y798 = n7890;
  assign y799 = n7896;
  assign y800 = n7902;
  assign y801 = n7908;
  assign y802 = n7914;
  assign y803 = n7920;
  assign y804 = n7926;
  assign y805 = n7932;
  assign y806 = n7938;
  assign y807 = n7944;
  assign y808 = n7950;
  assign y809 = n7956;
  assign y810 = n7962;
  assign y811 = n7968;
  assign y812 = n7974;
  assign y813 = n7980;
  assign y814 = n7986;
  assign y815 = n7992;
  assign y816 = ~n8002;
  assign y817 = n8008;
  assign y818 = n8014;
  assign y819 = n8020;
  assign y820 = ~n8072;
  assign y821 = ~n8118;
  assign y822 = n8124;
  assign y823 = ~n8172;
  assign y824 = ~n8227;
  assign y825 = ~n8280;
  assign y826 = n8286;
  assign y827 = ~n8320;
  assign y828 = ~n8355;
  assign y829 = ~n8408;
  assign y830 = ~n8454;
  assign y831 = ~n8508;
  assign y832 = ~n8556;
  assign y833 = ~n8609;
  assign y834 = ~n8649;
  assign y835 = ~n8682;
  assign y836 = ~n8729;
  assign y837 = n8735;
  assign y838 = n8741;
  assign y839 = ~n8776;
  assign y840 = n1478;
  assign y841 = n8783;
  assign y842 = ~n8831;
  assign y843 = n8837;
  assign y844 = n8843;
  assign y845 = n8849;
  assign y846 = ~n8899;
  assign y847 = n8905;
  assign y848 = n8911;
  assign y849 = ~n8954;
  assign y850 = n8960;
  assign y851 = n8966;
  assign y852 = n8972;
  assign y853 = n8978;
  assign y854 = n8984;
  assign y855 = n8990;
  assign y856 = n8996;
  assign y857 = n9002;
  assign y858 = n9008;
  assign y859 = n9014;
  assign y860 = n9020;
  assign y861 = n9026;
  assign y862 = n9032;
  assign y863 = n9038;
  assign y864 = ~n9077;
  assign y865 = ~n9123;
  assign y866 = n9129;
  assign y867 = n9135;
  assign y868 = ~n9174;
  assign y869 = ~n9213;
  assign y870 = ~n9252;
  assign y871 = ~n9307;
  assign y872 = n9313;
  assign y873 = ~n9352;
  assign y874 = ~n9404;
  assign y875 = ~n9443;
  assign y876 = ~n9497;
  assign y877 = ~n9552;
  assign y878 = n9575;
  assign y879 = ~n9623;
  assign y880 = n9629;
  assign y881 = n9635;
  assign y882 = n9641;
  assign y883 = n9647;
  assign y884 = n9653;
  assign y885 = n9659;
  assign y886 = n9665;
  assign y887 = n9671;
  assign y888 = n9675;
  assign y889 = n9681;
  assign y890 = ~n9727;
  assign y891 = n9733;
  assign y892 = n9739;
  assign y893 = n9745;
  assign y894 = n9751;
  assign y895 = n9757;
  assign y896 = ~n9764;
  assign y897 = n7636;
  assign y898 = ~n9770;
  assign y899 = ~n9776;
  assign y900 = ~n9782;
  assign y901 = ~n9788;
  assign y902 = ~n9794;
  assign y903 = ~n9800;
  assign y904 = n9803;
  assign y905 = ~n9809;
  assign y906 = ~n9815;
  assign y907 = ~n9821;
  assign y908 = ~n9827;
  assign y909 = ~n9833;
  assign y910 = ~n9839;
  assign y911 = ~n9845;
  assign y912 = ~n9851;
  assign y913 = ~n9857;
  assign y914 = ~n9863;
  assign y915 = ~n9869;
  assign y916 = ~n9875;
  assign y917 = ~n9881;
  assign y918 = ~n9887;
  assign y919 = ~n9893;
  assign y920 = ~n9899;
  assign y921 = ~n9905;
  assign y922 = n9915;
  assign y923 = ~n9921;
  assign y924 = ~n9927;
  assign y925 = ~n9933;
  assign y926 = n9935;
  assign y927 = ~n9941;
  assign y928 = n9945;
  assign y929 = ~n9951;
  assign y930 = n9953;
  assign y931 = ~n9959;
  assign y932 = n9963;
  assign y933 = ~n9969;
  assign y934 = ~n9975;
  assign y935 = n9983;
  assign y936 = ~n9984;
  assign y937 = ~n9985;
  assign y938 = n9988;
  assign y939 = ~n9990;
  assign y940 = n9993;
  assign y941 = n9996;
  assign y942 = n9999;
  assign y943 = ~n10002;
  assign y944 = n10005;
  assign y945 = n10008;
  assign y946 = n10011;
  assign y947 = n10014;
  assign y948 = n10017;
  assign y949 = n10020;
  assign y950 = n2390;
  assign y951 = n10024;
  assign y952 = n10027;
  assign y953 = ~n10034;
  assign y954 = n7788;
  assign y955 = n10037;
  assign y956 = ~n10040;
  assign y957 = n10043;
  assign y958 = n10046;
  assign y959 = n10047;
  assign y960 = ~n10050;
  assign y961 = n10053;
  assign y962 = ~n10054;
  assign y963 = n9913;
  assign y964 = n10057;
  assign y965 = n10060;
  assign y966 = ~n10063;
  assign y967 = n10066;
  assign y968 = n10069;
  assign y969 = ~n10072;
  assign y970 = n10075;
  assign y971 = ~n10078;
  assign y972 = n10081;
  assign y973 = n10084;
  assign y974 = ~n10085;
  assign y975 = ~n10086;
  assign y976 = ~n10087;
  assign y977 = ~n10089;
  assign y978 = n9574;
  assign y979 = n10090;
  assign y980 = n8777;
  assign y981 = n10094;
  assign y982 = ~n10105;
  assign y983 = ~n10115;
  assign y984 = ~n10125;
  assign y985 = ~n10135;
  assign y986 = ~n10139;
  assign y987 = ~n10140;
  assign y988 = n9758;
  assign y989 = n10143;
  assign y990 = n10146;
  assign y991 = n10147;
  assign y992 = ~n10149;
  assign y993 = n10152;
  assign y994 = n10155;
  assign y995 = n10158;
  assign y996 = n10161;
  assign y997 = n2959;
  assign y998 = n10164;
  assign y999 = n10167;
  assign y1000 = n10170;
  assign y1001 = n10173;
  assign y1002 = n10176;
  assign y1003 = n10179;
  assign y1004 = n10182;
  assign y1005 = n10185;
  assign y1006 = n10188;
  assign y1007 = n10191;
  assign y1008 = n10194;
  assign y1009 = n10197;
  assign y1010 = n10200;
  assign y1011 = n10203;
  assign y1012 = n10206;
  assign y1013 = n10209;
  assign y1014 = n10212;
  assign y1015 = n10215;
  assign y1016 = n10218;
  assign y1017 = n10221;
  assign y1018 = n10224;
  assign y1019 = n10227;
  assign y1020 = n10230;
  assign y1021 = n10233;
  assign y1022 = n10236;
  assign y1023 = n10239;
  assign y1024 = n10242;
  assign y1025 = n10245;
  assign y1026 = n10248;
  assign y1027 = n10251;
  assign y1028 = n10254;
  assign y1029 = n10257;
  assign y1030 = n10260;
  assign y1031 = n10263;
  assign y1032 = n10266;
  assign y1033 = n10269;
  assign y1034 = n10272;
  assign y1035 = n10275;
  assign y1036 = n10278;
  assign y1037 = n10281;
  assign y1038 = ~n1571;
  assign y1039 = ~n10284;
  assign y1040 = ~n10287;
  assign y1041 = ~n10290;
  assign y1042 = ~n10293;
  assign y1043 = ~n10296;
  assign y1044 = ~n10299;
  assign y1045 = ~n10302;
  assign y1046 = ~n10305;
  assign y1047 = ~n10308;
  assign y1048 = ~n10311;
  assign y1049 = ~n5523;
  assign y1050 = ~n10314;
  assign y1051 = ~n10317;
  assign y1052 = ~n10320;
  assign y1053 = x67;
  assign y1054 = ~n10323;
  assign y1055 = ~n10326;
  assign y1056 = ~n10329;
  assign y1057 = ~n2331;
  assign y1058 = ~n10332;
  assign y1059 = ~n10335;
  assign y1060 = ~n10338;
  assign y1061 = ~n10341;
  assign y1062 = ~n10344;
  assign y1063 = n10352;
  assign y1064 = ~n10355;
  assign y1065 = ~n10358;
  assign y1066 = ~n10361;
  assign y1067 = ~n10364;
  assign y1068 = ~n10367;
  assign y1069 = ~n10370;
  assign y1070 = ~n10371;
  assign y1071 = ~n10374;
  assign y1072 = ~n10377;
  assign y1073 = ~n10380;
  assign y1074 = ~n10383;
  assign y1075 = ~n10386;
  assign y1076 = n10389;
  assign y1077 = n10392;
  assign y1078 = n10395;
  assign y1079 = n10398;
  assign y1080 = n10399;
  assign y1081 = n10402;
  assign y1082 = n10405;
  assign y1083 = n10408;
  assign y1084 = n10411;
  assign y1085 = n10414;
  assign y1086 = n10417;
  assign y1087 = n10420;
  assign y1088 = n10422;
  assign y1089 = n10425;
  assign y1090 = n10428;
  assign y1091 = n10431;
  assign y1092 = n10434;
  assign y1093 = n10437;
  assign y1094 = n10440;
  assign y1095 = n10443;
  assign y1096 = n10446;
  assign y1097 = n10449;
  assign y1098 = n10452;
  assign y1099 = n10455;
  assign y1100 = n10458;
  assign y1101 = ~n2353;
  assign y1102 = n10459;
  assign y1103 = n10463;
  assign y1104 = n10464;
  assign y1105 = ~n10467;
  assign y1106 = n10468;
  assign y1107 = n2479;
  assign y1108 = x1134;
  assign y1109 = x964;
  assign y1110 = ~x954;
  assign y1111 = x965;
  assign y1112 = ~n10470;
  assign y1113 = x991;
  assign y1114 = x985;
  assign y1115 = n10471;
  assign y1116 = n10472;
  assign y1117 = x1014;
  assign y1118 = n10473;
  assign y1119 = x1029;
  assign y1120 = x1004;
  assign y1121 = x1007;
  assign y1122 = n10474;
  assign y1123 = x1135;
  assign y1124 = n10475;
  assign y1125 = n10476;
  assign y1126 = n10477;
  assign y1127 = n10478;
  assign y1128 = n10479;
  assign y1129 = n10480;
  assign y1130 = ~x278;
  assign y1131 = n10481;
  assign y1132 = n10482;
  assign y1133 = ~n10483;
  assign y1134 = x1064;
  assign y1135 = n10484;
  assign y1136 = x299;
  assign y1137 = ~n10485;
  assign y1138 = x1075;
  assign y1139 = x1052;
  assign y1140 = x771;
  assign y1141 = x765;
  assign y1142 = x605;
  assign y1143 = x601;
  assign y1144 = x278;
  assign y1145 = x279;
  assign y1146 = ~x915;
  assign y1147 = ~x825;
  assign y1148 = ~x826;
  assign y1149 = ~x913;
  assign y1150 = ~x894;
  assign y1151 = ~x905;
  assign y1152 = x1095;
  assign y1153 = ~x890;
  assign y1154 = x1094;
  assign y1155 = ~x906;
  assign y1156 = ~x896;
  assign y1157 = ~x909;
  assign y1158 = ~x911;
  assign y1159 = ~x908;
  assign y1160 = ~x891;
  assign y1161 = ~x902;
  assign y1162 = ~x903;
  assign y1163 = ~x883;
  assign y1164 = ~x888;
  assign y1165 = ~x919;
  assign y1166 = ~x886;
  assign y1167 = ~x912;
  assign y1168 = ~x895;
  assign y1169 = ~x916;
  assign y1170 = ~x889;
  assign y1171 = ~x900;
  assign y1172 = ~x885;
  assign y1173 = ~x904;
  assign y1174 = ~x899;
  assign y1175 = ~x918;
  assign y1176 = ~x898;
  assign y1177 = ~x917;
  assign y1178 = ~x827;
  assign y1179 = ~x887;
  assign y1180 = ~x884;
  assign y1181 = ~x910;
  assign y1182 = ~x828;
  assign y1183 = ~x892;
  assign y1184 = x1187;
  assign y1185 = x1172;
  assign y1186 = x1170;
  assign y1187 = x1138;
  assign y1188 = x1177;
  assign y1189 = x1178;
  assign y1190 = x863;
  assign y1191 = x1203;
  assign y1192 = x1185;
  assign y1193 = x1171;
  assign y1194 = x1192;
  assign y1195 = x1137;
  assign y1196 = x1186;
  assign y1197 = x1165;
  assign y1198 = x1164;
  assign y1199 = x1098;
  assign y1200 = x1183;
  assign y1201 = x230;
  assign y1202 = x1169;
  assign y1203 = x1136;
  assign y1204 = x1181;
  assign y1205 = x849;
  assign y1206 = x1193;
  assign y1207 = x1182;
  assign y1208 = x1168;
  assign y1209 = x1175;
  assign y1210 = x1191;
  assign y1211 = x1099;
  assign y1212 = x1174;
  assign y1213 = x1179;
  assign y1214 = x1202;
  assign y1215 = x1176;
  assign y1216 = x1173;
  assign y1217 = x1201;
  assign y1218 = x1167;
  assign y1219 = x840;
  assign y1220 = x1189;
  assign y1221 = x1195;
  assign y1222 = x864;
  assign y1223 = x1190;
  assign y1224 = x1188;
  assign y1225 = x1180;
  assign y1226 = x1194;
  assign y1227 = x1097;
  assign y1228 = x1166;
  assign y1229 = x1200;
  assign y1230 = x1184;
endmodule