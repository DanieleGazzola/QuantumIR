module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869;
  assign n25 = ~x0 & ~x1;
  assign n26 = ~x2 & n25;
  assign n27 = ~x3 & n26;
  assign n28 = ~x4 & n27;
  assign n34 = ~x5 & n28;
  assign n35 = ~x6 & ~x7;
  assign n36 = n34 & n35;
  assign n37 = ~x8 & n36;
  assign n38 = ~x9 & n37;
  assign n39 = ~x10 & n38;
  assign n40 = ~x11 & n39;
  assign n41 = ~x12 & ~x13;
  assign n42 = ~x14 & n41;
  assign n43 = n40 & n42;
  assign n44 = ~x22 & ~n43;
  assign n45 = n44 ^ x15;
  assign n46 = ~x15 & n43;
  assign n47 = ~x22 & ~n46;
  assign n48 = ~x18 & ~x19;
  assign n49 = ~x16 & ~x17;
  assign n50 = n48 & n49;
  assign n51 = ~n47 & n50;
  assign n52 = ~x22 & ~n51;
  assign n53 = n52 ^ x20;
  assign n54 = x22 ^ x21;
  assign n55 = n53 & n54;
  assign n56 = ~n45 & n55;
  assign n57 = x21 ^ x20;
  assign n58 = n52 ^ x21;
  assign n59 = n57 & n58;
  assign n60 = n45 & n59;
  assign n61 = ~n56 & ~n60;
  assign n62 = n46 ^ x16;
  assign n63 = x17 & ~n62;
  assign n64 = x19 & ~x22;
  assign n65 = ~x18 & n64;
  assign n66 = n63 & n65;
  assign n67 = x16 & ~x17;
  assign n68 = x18 & ~x19;
  assign n69 = x22 & n68;
  assign n70 = n67 & n69;
  assign n71 = ~n66 & ~n70;
  assign n72 = ~x22 & n68;
  assign n73 = x17 ^ x16;
  assign n74 = n46 ^ x17;
  assign n75 = n73 & ~n74;
  assign n76 = n72 & n75;
  assign n77 = ~x18 & x19;
  assign n78 = x22 & n77;
  assign n79 = ~x16 & x17;
  assign n80 = n78 & n79;
  assign n81 = ~n76 & ~n80;
  assign n82 = n71 & n81;
  assign n83 = ~n45 & n81;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~n61 & n84;
  assign n86 = ~n45 & n59;
  assign n171 = n45 & ~n54;
  assign n172 = n53 & n171;
  assign n89 = x18 & x19;
  assign n132 = ~x22 & n89;
  assign n268 = n63 & n132;
  assign n134 = x22 & n48;
  assign n269 = n67 & n134;
  assign n270 = ~n268 & ~n269;
  assign n319 = n172 & ~n270;
  assign n320 = ~n86 & ~n319;
  assign n321 = ~n85 & n320;
  assign n118 = n65 & n75;
  assign n119 = n69 & n79;
  assign n120 = ~n118 & ~n119;
  assign n322 = n83 & n120;
  assign n323 = ~n321 & ~n322;
  assign n94 = n54 & ~n57;
  assign n184 = n45 & n94;
  assign n143 = n46 ^ x18;
  assign n144 = n143 ^ x22;
  assign n145 = n49 ^ n46;
  assign n146 = n145 ^ n49;
  assign n96 = x16 & x17;
  assign n147 = n96 ^ n49;
  assign n148 = ~n146 & n147;
  assign n149 = n148 ^ n49;
  assign n150 = n149 ^ n143;
  assign n151 = n144 & ~n150;
  assign n152 = n151 ^ n148;
  assign n153 = n152 ^ n49;
  assign n154 = n153 ^ x22;
  assign n155 = ~n143 & ~n154;
  assign n156 = n155 ^ n143;
  assign n217 = n49 & n89;
  assign n218 = n156 & ~n217;
  assign n219 = ~n64 & ~n218;
  assign n248 = n184 & n219;
  assign n112 = ~x17 & ~n62;
  assign n133 = n112 & n132;
  assign n135 = n96 & n134;
  assign n136 = ~n133 & ~n135;
  assign n249 = n86 & ~n136;
  assign n250 = ~n248 & ~n249;
  assign n87 = ~x22 & n48;
  assign n88 = n75 & n87;
  assign n90 = x22 & n89;
  assign n91 = n79 & n90;
  assign n92 = ~n88 & ~n91;
  assign n324 = n61 & ~n92;
  assign n325 = n250 & ~n324;
  assign n139 = n75 & n132;
  assign n140 = n79 & n134;
  assign n141 = ~n139 & ~n140;
  assign n326 = ~n141 & n184;
  assign n106 = n45 & n55;
  assign n327 = n106 & ~n270;
  assign n328 = ~n326 & ~n327;
  assign n329 = n325 & n328;
  assign n330 = ~n323 & n329;
  assign n331 = ~n56 & n330;
  assign n97 = ~n46 & n96;
  assign n162 = n97 & n132;
  assign n163 = ~n51 & ~n162;
  assign n164 = n65 & n112;
  assign n165 = n69 & n96;
  assign n166 = ~n164 & ~n165;
  assign n167 = n163 & n166;
  assign n332 = n167 & ~n172;
  assign n333 = ~n331 & ~n332;
  assign n157 = x19 & ~n156;
  assign n158 = n49 & n69;
  assign n159 = ~n157 & ~n158;
  assign n334 = n92 & n159;
  assign n335 = n163 & n270;
  assign n336 = n136 & n141;
  assign n337 = n335 & n336;
  assign n338 = n59 & n337;
  assign n95 = ~n45 & n94;
  assign n176 = n87 & n112;
  assign n177 = n90 & n96;
  assign n178 = ~n176 & ~n177;
  assign n287 = n63 & n87;
  assign n288 = n67 & n90;
  assign n289 = ~n287 & ~n288;
  assign n339 = n178 & n289;
  assign n340 = n92 & n339;
  assign n341 = n95 & n340;
  assign n342 = ~n338 & ~n341;
  assign n343 = n334 & n342;
  assign n109 = n53 & ~n54;
  assign n110 = ~n45 & n109;
  assign n344 = n71 & ~n110;
  assign n345 = ~n343 & ~n344;
  assign n113 = n72 & n112;
  assign n114 = n78 & n96;
  assign n115 = ~n113 & ~n114;
  assign n346 = n115 & n159;
  assign n347 = n141 & n346;
  assign n348 = n172 & ~n347;
  assign n349 = n92 & n166;
  assign n350 = ~n86 & n349;
  assign n351 = n71 & ~n184;
  assign n352 = n120 & n351;
  assign n353 = ~n350 & ~n352;
  assign n354 = ~n348 & ~n353;
  assign n111 = ~n81 & n110;
  assign n116 = n110 & ~n115;
  assign n117 = ~n111 & ~n116;
  assign n355 = n110 & ~n136;
  assign n356 = n117 & ~n355;
  assign n357 = n354 & n356;
  assign n358 = ~n345 & n357;
  assign n359 = ~n333 & n358;
  assign n436 = n86 & ~n270;
  assign n818 = n71 & ~n436;
  assign n819 = ~n86 & ~n95;
  assign n820 = ~n818 & ~n819;
  assign n142 = n56 & ~n141;
  assign n821 = ~n142 & ~n248;
  assign n822 = ~n820 & n821;
  assign n93 = n86 & ~n92;
  assign n823 = ~n55 & ~n60;
  assign n824 = ~n115 & ~n823;
  assign n825 = ~n93 & ~n824;
  assign n681 = n86 & n219;
  assign n647 = n184 & ~n270;
  assign n655 = n136 & n289;
  assign n826 = n95 & ~n655;
  assign n827 = ~n647 & ~n826;
  assign n828 = n141 & n178;
  assign n829 = n106 & ~n828;
  assign n830 = n827 & ~n829;
  assign n831 = ~n681 & n830;
  assign n832 = n825 & n831;
  assign n833 = n822 & n832;
  assign n834 = ~n86 & n833;
  assign n667 = ~n86 & ~n184;
  assign n668 = ~n159 & ~n667;
  assign n835 = ~n184 & ~n219;
  assign n836 = ~n668 & n835;
  assign n837 = ~n834 & ~n836;
  assign n444 = n60 & ~n270;
  assign n121 = n63 & n72;
  assign n122 = n67 & n78;
  assign n123 = ~n121 & ~n122;
  assign n185 = ~n123 & n184;
  assign n374 = n95 & ~n159;
  assign n1054 = ~n185 & ~n374;
  assign n1055 = ~n444 & n1054;
  assign n173 = ~n81 & n172;
  assign n174 = ~n81 & n95;
  assign n175 = ~n173 & ~n174;
  assign n547 = ~n60 & n163;
  assign n838 = n81 & n92;
  assign n839 = ~n172 & n838;
  assign n840 = ~n547 & ~n839;
  assign n2024 = n175 & ~n840;
  assign n2025 = n1055 & n2024;
  assign n98 = n72 & n97;
  assign n99 = n49 & n77;
  assign n100 = ~n47 & n99;
  assign n101 = ~n98 & ~n100;
  assign n472 = ~n101 & n110;
  assign n403 = n95 & ~n289;
  assign n1049 = n86 & ~n163;
  assign n1268 = ~n403 & ~n1049;
  assign n1269 = ~n472 & n1268;
  assign n687 = n106 & ~n115;
  assign n124 = n120 & n123;
  assign n125 = n110 & ~n124;
  assign n198 = n56 & ~n178;
  assign n2026 = ~n125 & ~n198;
  assign n2027 = ~n687 & n2026;
  assign n2028 = n1269 & n2027;
  assign n2029 = n2025 & n2028;
  assign n2030 = ~n837 & n2029;
  assign n408 = n115 & n178;
  assign n409 = n110 & ~n408;
  assign n410 = ~n166 & n184;
  assign n411 = ~n409 & ~n410;
  assign n256 = n120 & n166;
  assign n412 = n106 & ~n256;
  assign n413 = n411 & ~n412;
  assign n294 = n86 & ~n178;
  assign n414 = n110 & ~n163;
  assign n415 = ~n294 & ~n414;
  assign n203 = n45 & ~n141;
  assign n204 = n59 & n203;
  assign n207 = ~n45 & ~n123;
  assign n416 = n55 & n207;
  assign n417 = ~n204 & ~n416;
  assign n290 = ~n219 & n289;
  assign n418 = n172 & ~n290;
  assign n419 = n417 & ~n418;
  assign n420 = n415 & n419;
  assign n421 = n413 & n420;
  assign n260 = ~n163 & n184;
  assign n510 = n95 & ~n141;
  assign n360 = n106 & ~n166;
  assign n362 = n56 & ~n81;
  assign n3454 = ~n360 & ~n362;
  assign n3455 = ~n510 & n3454;
  assign n3786 = ~n260 & n3455;
  assign n105 = n56 & ~n71;
  assign n1980 = ~n105 & ~n326;
  assign n208 = n59 & n207;
  assign n659 = n60 & ~n289;
  assign n2237 = ~n208 & ~n659;
  assign n3787 = ~n93 & n2237;
  assign n3788 = n1980 & n3787;
  assign n3789 = n3786 & n3788;
  assign n507 = ~n136 & n184;
  assign n199 = ~n81 & n86;
  assign n314 = ~n120 & n172;
  assign n628 = n56 & ~n136;
  assign n1270 = ~n314 & ~n628;
  assign n1271 = ~n199 & n1270;
  assign n1994 = ~n507 & n1271;
  assign n235 = n60 & ~n120;
  assign n3065 = ~n110 & n141;
  assign n3066 = n71 & ~n106;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = ~n235 & ~n3067;
  assign n255 = n60 & ~n178;
  assign n371 = n60 & ~n163;
  assign n3069 = ~n255 & ~n371;
  assign n3070 = n3068 & n3069;
  assign n3790 = n1994 & n3070;
  assign n3791 = n3789 & n3790;
  assign n3792 = n421 & n3791;
  assign n3793 = n2030 & n3792;
  assign n3794 = n359 & n3793;
  assign n2321 = x22 ^ x2;
  assign n2322 = ~x1 & x2;
  assign n2323 = n2321 & ~n2322;
  assign n3118 = x2 ^ x1;
  assign n3267 = x0 & ~n3118;
  assign n422 = n92 & ~n219;
  assign n423 = n45 & ~n422;
  assign n424 = n340 & ~n423;
  assign n425 = n94 & ~n424;
  assign n426 = n56 & ~n163;
  assign n427 = n71 & n159;
  assign n428 = n59 & ~n427;
  assign n429 = ~n426 & ~n428;
  assign n430 = ~n425 & n429;
  assign n548 = ~n106 & n427;
  assign n549 = ~n547 & ~n548;
  assign n550 = n430 & ~n549;
  assign n2389 = n159 & n336;
  assign n3100 = n270 & n2389;
  assign n3101 = n55 & ~n3100;
  assign n3102 = n550 & ~n3101;
  assign n285 = n109 & ~n136;
  assign n286 = ~n173 & ~n285;
  assign n291 = n60 & ~n290;
  assign n292 = n286 & ~n291;
  assign n293 = n117 & n292;
  assign n295 = n92 & ~n109;
  assign n296 = ~n294 & n295;
  assign n297 = ~n59 & ~n219;
  assign n298 = ~n115 & n172;
  assign n299 = n297 & ~n298;
  assign n300 = ~n296 & ~n299;
  assign n301 = n86 & ~n290;
  assign n302 = ~n300 & ~n301;
  assign n303 = n293 & n302;
  assign n535 = n115 & n289;
  assign n536 = ~n423 & n535;
  assign n537 = n55 & ~n536;
  assign n538 = ~n198 & ~n537;
  assign n3103 = n120 & n427;
  assign n3104 = ~n59 & ~n110;
  assign n3105 = ~n3103 & ~n3104;
  assign n252 = ~n123 & n172;
  assign n711 = ~n159 & n172;
  assign n3106 = ~n252 & ~n711;
  assign n3107 = ~n3105 & n3106;
  assign n232 = n60 & ~n166;
  assign n233 = ~n71 & n172;
  assign n234 = ~n232 & ~n233;
  assign n845 = n86 & ~n166;
  assign n3108 = n56 & ~n422;
  assign n3109 = ~n845 & ~n3108;
  assign n3110 = n234 & n3109;
  assign n3111 = n3107 & n3110;
  assign n3112 = n538 & n3111;
  assign n3113 = n303 & n3112;
  assign n3114 = n3102 & n3113;
  assign n539 = n56 & n219;
  assign n1977 = ~n436 & ~n539;
  assign n622 = n86 & ~n289;
  assign n1978 = ~n622 & ~n687;
  assign n1979 = n1977 & n1978;
  assign n654 = n56 & ~n289;
  assign n872 = ~n371 & ~n654;
  assign n1981 = n872 & n1980;
  assign n1982 = n1979 & n1981;
  assign n304 = n159 & n166;
  assign n305 = ~n59 & n304;
  assign n306 = n101 & n123;
  assign n307 = ~n109 & n306;
  assign n308 = ~n305 & ~n307;
  assign n2087 = n94 & ~n270;
  assign n2088 = n163 & ~n2087;
  assign n887 = n56 & ~n115;
  assign n3046 = n109 & ~n289;
  assign n3047 = ~n887 & ~n3046;
  assign n3048 = n2088 & n3047;
  assign n3049 = ~n308 & n3048;
  assign n315 = ~n255 & ~n314;
  assign n214 = n106 & ~n120;
  assign n707 = ~n214 & ~n507;
  assign n3050 = n315 & n707;
  assign n3051 = n3049 & n3050;
  assign n227 = ~n92 & n110;
  assign n488 = n95 & ~n136;
  assign n642 = ~n444 & ~n488;
  assign n3052 = ~n227 & n642;
  assign n2249 = ~n374 & ~n510;
  assign n1901 = n106 & n219;
  assign n3053 = ~n252 & ~n1901;
  assign n3054 = n2249 & n3053;
  assign n3055 = n3052 & n3054;
  assign n3056 = n3051 & n3055;
  assign n3057 = n1982 & n3056;
  assign n474 = n106 & ~n178;
  assign n1083 = ~n360 & ~n474;
  assign n131 = ~n71 & n106;
  assign n2085 = n56 & ~n256;
  assign n2086 = ~n131 & ~n2085;
  assign n3058 = n1083 & n2086;
  assign n367 = n110 & ~n270;
  assign n3059 = ~n367 & ~n681;
  assign n3060 = n3058 & n3059;
  assign n3061 = n293 & n3060;
  assign n3062 = n550 & n3061;
  assign n3063 = n3057 & n3062;
  assign n1272 = n1269 & n1271;
  assign n451 = n45 & n53;
  assign n452 = ~n289 & n451;
  assign n453 = n54 & n452;
  assign n454 = n71 & n136;
  assign n455 = ~n219 & n454;
  assign n456 = n86 & ~n455;
  assign n457 = ~n453 & ~n456;
  assign n179 = n95 & ~n178;
  assign n506 = n106 & ~n136;
  assign n1273 = ~n506 & ~n622;
  assign n1274 = ~n179 & n1273;
  assign n1275 = n457 & n1274;
  assign n1276 = n1272 & n1275;
  assign n274 = n86 & ~n101;
  assign n1063 = n172 & ~n335;
  assign n1064 = ~n647 & ~n1063;
  assign n1277 = n92 & n1064;
  assign n1278 = n171 & ~n1277;
  assign n1279 = ~n274 & ~n1278;
  assign n1280 = n1276 & n1279;
  assign n278 = ~n71 & n95;
  assign n464 = n56 & ~n101;
  assign n2076 = ~n278 & ~n464;
  assign n379 = n106 & ~n123;
  assign n459 = ~n81 & n184;
  assign n2077 = ~n379 & ~n459;
  assign n2078 = n2076 & n2077;
  assign n2079 = ~n539 & ~n845;
  assign n2080 = ~n668 & n2079;
  assign n2081 = n2078 & n2080;
  assign n205 = ~n71 & n184;
  assign n727 = n109 & n207;
  assign n2082 = ~n205 & ~n727;
  assign n2083 = ~n214 & n2082;
  assign n2084 = n2081 & n2083;
  assign n183 = n86 & ~n115;
  assign n1284 = ~n183 & ~n474;
  assign n551 = n115 & n123;
  assign n2386 = n172 & ~n551;
  assign n2387 = ~n174 & ~n2386;
  assign n2388 = n1284 & n2387;
  assign n2390 = n290 & n2389;
  assign n2391 = n110 & ~n2390;
  assign n2392 = n2388 & ~n2391;
  assign n2393 = n2084 & n2392;
  assign n180 = n86 & ~n141;
  assign n241 = n110 & ~n141;
  assign n433 = ~n180 & ~n241;
  assign n434 = ~n120 & n184;
  assign n435 = n433 & ~n434;
  assign n437 = ~n255 & ~n436;
  assign n438 = ~n178 & n184;
  assign n439 = ~n82 & n172;
  assign n440 = ~n438 & ~n439;
  assign n441 = n437 & n440;
  assign n442 = n435 & n441;
  assign n107 = ~n92 & n106;
  assign n108 = ~n105 & ~n107;
  assign n682 = n86 & ~n120;
  assign n1020 = n55 & ~n270;
  assign n1021 = ~n682 & ~n1020;
  assign n1022 = n108 & n1021;
  assign n1924 = ~n185 & ~n208;
  assign n2394 = ~n290 & ~n667;
  assign n363 = n172 & ~n178;
  assign n397 = n95 & ~n166;
  assign n501 = n95 & ~n120;
  assign n2395 = ~n397 & ~n501;
  assign n2396 = ~n363 & n2395;
  assign n2397 = ~n887 & n2396;
  assign n2398 = ~n2394 & n2397;
  assign n2399 = n1924 & n2398;
  assign n2400 = n1022 & n2399;
  assign n2401 = n442 & n2400;
  assign n2402 = n2393 & n2401;
  assign n2403 = n1280 & n2402;
  assign n726 = ~n326 & ~n549;
  assign n251 = ~n71 & n110;
  assign n368 = ~n45 & n53;
  assign n1902 = ~n109 & ~n368;
  assign n1903 = ~n163 & ~n1902;
  assign n1904 = ~n1901 & ~n1903;
  assign n1905 = ~n251 & n1904;
  assign n1906 = n726 & n1905;
  assign n904 = n178 & ~n219;
  assign n905 = n110 & ~n904;
  assign n906 = ~n227 & ~n905;
  assign n1907 = n906 & n1021;
  assign n386 = n101 & ~n184;
  assign n673 = ~n106 & n120;
  assign n674 = ~n386 & ~n673;
  assign n1908 = ~n410 & ~n674;
  assign n1909 = n1907 & n1908;
  assign n1910 = n1906 & n1909;
  assign n479 = n56 & ~n92;
  assign n669 = ~n274 & ~n479;
  assign n126 = n60 & ~n92;
  assign n1911 = ~n126 & ~n131;
  assign n1912 = n669 & n1911;
  assign n1913 = ~n453 & ~n501;
  assign n1914 = n1912 & n1913;
  assign n1915 = n1910 & n1914;
  assign n398 = ~n101 & n172;
  assign n1916 = ~n241 & ~n398;
  assign n1917 = ~n360 & n1916;
  assign n1918 = ~n179 & ~n845;
  assign n1919 = ~n668 & n1918;
  assign n1920 = n1917 & n1919;
  assign n1921 = n833 & n1920;
  assign n1922 = n1915 & n1921;
  assign n390 = ~n45 & ~n120;
  assign n1012 = n109 & n390;
  assign n1923 = ~n198 & ~n1012;
  assign n1925 = n71 & n166;
  assign n1926 = n56 & ~n1925;
  assign n1927 = n1924 & ~n1926;
  assign n1928 = n1923 & n1927;
  assign n1283 = ~n444 & ~n510;
  assign n491 = n60 & n219;
  assign n1929 = ~n379 & ~n491;
  assign n1930 = n1283 & n1929;
  assign n1931 = n1928 & n1930;
  assign n688 = ~n438 & ~n687;
  assign n220 = ~n166 & n171;
  assign n689 = ~n55 & n115;
  assign n690 = ~n94 & n136;
  assign n691 = ~n45 & ~n690;
  assign n692 = ~n689 & n691;
  assign n693 = ~n220 & ~n692;
  assign n694 = n688 & n693;
  assign n1932 = n117 & ~n235;
  assign n267 = n60 & ~n101;
  assign n445 = n110 & ~n289;
  assign n650 = ~n267 & ~n445;
  assign n554 = ~n101 & n184;
  assign n626 = n123 & n136;
  assign n1933 = n172 & ~n626;
  assign n1934 = ~n554 & ~n1933;
  assign n1935 = n650 & n1934;
  assign n1936 = n1932 & n1935;
  assign n1937 = n694 & n1936;
  assign n1938 = n1931 & n1937;
  assign n1939 = n1922 & n1938;
  assign n309 = n115 & n166;
  assign n310 = n81 & n309;
  assign n311 = n59 & ~n310;
  assign n312 = ~n235 & ~n311;
  assign n313 = ~n308 & n312;
  assign n316 = ~n109 & n315;
  assign n317 = n313 & n316;
  assign n318 = n303 & n317;
  assign n534 = n59 & n318;
  assign n540 = n86 & ~n337;
  assign n541 = ~n479 & ~n540;
  assign n512 = n81 & n178;
  assign n542 = n106 & ~n512;
  assign n543 = n541 & ~n542;
  assign n544 = ~n539 & n543;
  assign n545 = n538 & n544;
  assign n546 = ~n534 & n545;
  assign n552 = n81 & n551;
  assign n553 = n94 & ~n552;
  assign n473 = n95 & n219;
  assign n555 = ~n473 & ~n554;
  assign n556 = ~n553 & n555;
  assign n557 = n550 & n556;
  assign n558 = n546 & n557;
  assign n102 = n95 & ~n101;
  assign n361 = ~n102 & ~n360;
  assign n364 = ~n362 & ~n363;
  assign n365 = n361 & n364;
  assign n366 = n359 & n365;
  assign n369 = ~n101 & n368;
  assign n370 = ~n367 & ~n369;
  assign n372 = ~n205 & ~n371;
  assign n373 = n370 & n372;
  assign n375 = n60 & ~n159;
  assign n376 = ~n374 & ~n375;
  assign n377 = n250 & n376;
  assign n378 = n373 & n377;
  assign n380 = n109 & ~n167;
  assign n381 = ~n110 & ~n380;
  assign n382 = ~n379 & n381;
  assign n383 = ~n45 & n71;
  assign n384 = ~n382 & ~n383;
  assign n385 = ~n106 & n159;
  assign n387 = n163 & n386;
  assign n388 = ~n385 & ~n387;
  assign n389 = n109 & ~n124;
  assign n186 = ~n92 & n95;
  assign n391 = ~n186 & ~n390;
  assign n392 = ~n389 & n391;
  assign n393 = ~n388 & n392;
  assign n394 = ~n384 & n393;
  assign n395 = n378 & n394;
  assign n396 = n366 & n395;
  assign n137 = n60 & ~n136;
  assign n138 = ~n131 & ~n137;
  assign n399 = n110 & ~n166;
  assign n400 = ~n398 & ~n399;
  assign n401 = ~n397 & n400;
  assign n402 = n138 & n401;
  assign n404 = ~n110 & n163;
  assign n405 = ~n297 & ~n404;
  assign n406 = ~n403 & ~n405;
  assign n407 = n402 & n406;
  assign n431 = n421 & n430;
  assign n432 = n407 & n431;
  assign n443 = ~n136 & n172;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n443 & n446;
  assign n448 = n442 & n447;
  assign n449 = n432 & n448;
  assign n450 = n396 & n449;
  assign n103 = ~n93 & ~n102;
  assign n104 = ~n85 & n103;
  assign n458 = n104 & n457;
  assign n460 = n109 & ~n178;
  assign n461 = ~n45 & n460;
  assign n462 = ~n459 & ~n461;
  assign n463 = ~n416 & n462;
  assign n465 = n106 & ~n159;
  assign n466 = ~n464 & ~n465;
  assign n467 = n463 & n466;
  assign n468 = n458 & n467;
  assign n469 = n136 & n346;
  assign n470 = n60 & ~n469;
  assign n471 = ~n314 & ~n470;
  assign n475 = ~n473 & ~n474;
  assign n476 = ~n472 & n475;
  assign n477 = n471 & n476;
  assign n478 = n468 & n477;
  assign n127 = ~n125 & ~n126;
  assign n128 = n117 & n127;
  assign n129 = n108 & n128;
  assign n195 = n166 & ~n172;
  assign n196 = n92 & ~n184;
  assign n197 = ~n195 & ~n196;
  assign n480 = ~n445 & ~n479;
  assign n481 = ~n197 & n480;
  assign n482 = n166 & ~n184;
  assign n483 = ~n252 & n482;
  assign n484 = ~n109 & n120;
  assign n485 = ~n483 & ~n484;
  assign n486 = n481 & ~n485;
  assign n487 = n129 & n486;
  assign n489 = ~n397 & ~n488;
  assign n490 = ~n198 & n489;
  assign n492 = n56 & ~n334;
  assign n493 = ~n491 & ~n492;
  assign n494 = ~n101 & n451;
  assign n495 = ~n426 & ~n494;
  assign n496 = n493 & n495;
  assign n497 = n490 & n496;
  assign n498 = n487 & n497;
  assign n499 = n478 & n498;
  assign n500 = ~n71 & n109;
  assign n502 = ~n326 & ~n501;
  assign n503 = ~n500 & n502;
  assign n209 = ~n115 & n184;
  assign n504 = ~n179 & ~n209;
  assign n505 = n503 & n504;
  assign n508 = ~n438 & ~n507;
  assign n509 = ~n506 & n508;
  assign n511 = ~n227 & ~n510;
  assign n513 = n115 & n512;
  assign n514 = n172 & ~n513;
  assign n515 = n289 & ~n390;
  assign n516 = n59 & ~n515;
  assign n517 = ~n514 & ~n516;
  assign n518 = n511 & n517;
  assign n519 = n509 & n518;
  assign n520 = n505 & n519;
  assign n521 = n172 & ~n289;
  assign n522 = n110 & n219;
  assign n523 = ~n379 & ~n522;
  assign n524 = ~n521 & n523;
  assign n264 = n172 & n219;
  assign n525 = n106 & ~n163;
  assign n526 = ~n264 & ~n525;
  assign n277 = n95 & ~n115;
  assign n527 = ~n86 & ~n277;
  assign n528 = ~n346 & ~n527;
  assign n529 = n526 & ~n528;
  assign n530 = n524 & n529;
  assign n531 = n520 & n530;
  assign n532 = n499 & n531;
  assign n592 = ~n450 & ~n532;
  assign n593 = ~n558 & ~n592;
  assign n594 = ~x22 & ~n39;
  assign n595 = n594 ^ x11;
  assign n560 = ~x22 & ~n40;
  assign n579 = n560 ^ x12;
  assign n596 = n595 ^ n579;
  assign n597 = ~n318 & n596;
  assign n598 = ~n593 & ~n597;
  assign n571 = ~n55 & n558;
  assign n561 = x12 & ~x22;
  assign n562 = ~n560 & ~n561;
  assign n572 = n562 ^ x13;
  assign n563 = x13 & ~x22;
  assign n564 = n562 & ~n563;
  assign n565 = n564 ^ x14;
  assign n573 = n572 ^ n565;
  assign n574 = n546 & n573;
  assign n575 = n574 ^ n572;
  assign n576 = ~n571 & ~n575;
  assign n577 = ~n318 & n572;
  assign n578 = ~n576 & ~n577;
  assign n604 = n598 ^ n578;
  assign n533 = n532 ^ n450;
  assign n559 = n558 ^ n450;
  assign n566 = n565 ^ n450;
  assign n567 = n559 & n566;
  assign n568 = n567 ^ n450;
  assign n569 = ~n533 & ~n568;
  assign n570 = n569 ^ n558;
  assign n580 = ~n318 & ~n579;
  assign n581 = n571 & ~n580;
  assign n582 = n579 ^ n572;
  assign n583 = n582 ^ n579;
  assign n584 = n579 ^ n318;
  assign n585 = n584 ^ n579;
  assign n586 = n583 & n585;
  assign n587 = n586 ^ n579;
  assign n588 = n546 & ~n587;
  assign n589 = n588 ^ n579;
  assign n590 = ~n581 & n589;
  assign n605 = n570 & ~n590;
  assign n606 = ~n604 & n605;
  assign n792 = n318 & n604;
  assign n793 = ~n578 & n598;
  assign n794 = ~n595 & n793;
  assign n795 = ~n792 & ~n794;
  assign n796 = n590 & ~n795;
  assign n797 = ~n606 & ~n796;
  assign n599 = n572 & ~n598;
  assign n591 = n578 & ~n590;
  assign n600 = n599 ^ n591;
  assign n601 = n570 & n600;
  assign n602 = n601 ^ n591;
  assign n603 = ~n318 & n602;
  assign n607 = n578 & ~n598;
  assign n798 = ~n607 & ~n792;
  assign n799 = ~n570 & ~n798;
  assign n800 = ~n603 & ~n799;
  assign n801 = n797 & n800;
  assign n754 = n546 & ~n571;
  assign n755 = n579 & n754;
  assign n756 = n546 ^ n318;
  assign n757 = n595 & n756;
  assign n758 = n757 ^ n318;
  assign n759 = ~n755 & n758;
  assign n745 = n558 & n592;
  assign n746 = n450 & n532;
  assign n747 = ~n558 & n746;
  assign n748 = ~n745 & ~n747;
  assign n749 = n572 ^ n558;
  assign n750 = ~n748 & n749;
  assign n751 = n565 ^ n558;
  assign n752 = n533 & n751;
  assign n753 = ~n750 & ~n752;
  assign n760 = n759 ^ n753;
  assign n619 = ~x22 & ~n37;
  assign n620 = n619 ^ x9;
  assign n765 = ~n318 & n620;
  assign n761 = n579 ^ n558;
  assign n762 = ~n748 & ~n761;
  assign n763 = n533 & n749;
  assign n764 = ~n762 & ~n763;
  assign n766 = n765 ^ n764;
  assign n670 = ~n668 & n669;
  assign n671 = ~n205 & ~n474;
  assign n672 = n670 & n671;
  assign n675 = ~n403 & ~n674;
  assign n676 = n95 & ~n123;
  assign n677 = ~n105 & ~n676;
  assign n678 = ~n355 & n677;
  assign n679 = n675 & n678;
  assign n680 = n672 & n679;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~n199 & n683;
  assign n685 = n401 & n684;
  assign n686 = n680 & n685;
  assign n695 = ~n110 & ~n184;
  assign n696 = ~n335 & ~n695;
  assign n697 = ~n174 & ~n473;
  assign n698 = ~n654 & n697;
  assign n699 = ~n696 & n698;
  assign n160 = n56 & ~n159;
  assign n700 = ~n160 & ~n443;
  assign n701 = n699 & n700;
  assign n702 = n694 & n701;
  assign n703 = ~n436 & ~n659;
  assign n704 = n92 & ~n204;
  assign n705 = n703 & n704;
  assign n706 = n59 & ~n705;
  assign n708 = n159 & n270;
  assign n709 = n110 & ~n708;
  assign n710 = ~n105 & ~n709;
  assign n712 = ~n163 & n172;
  assign n713 = ~n711 & ~n712;
  assign n714 = n710 & n713;
  assign n715 = n707 & n714;
  assign n716 = ~n706 & n715;
  assign n717 = n702 & n716;
  assign n718 = n686 & n717;
  assign n719 = ~n95 & ~n110;
  assign n720 = ~n101 & ~n719;
  assign n721 = ~n92 & n184;
  assign n722 = n56 & ~n124;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~n720 & n723;
  assign n725 = ~n327 & n724;
  assign n638 = n166 & ~n219;
  assign n639 = n141 & n638;
  assign n640 = n106 & ~n639;
  assign n728 = ~n640 & ~n727;
  assign n729 = n726 & n728;
  assign n730 = n725 & n729;
  assign n731 = n60 & ~n551;
  assign n732 = ~n362 & ~n731;
  assign n733 = ~n186 & ~n647;
  assign n734 = n732 & n733;
  assign n735 = n730 & n734;
  assign n736 = n718 & n735;
  assign n623 = ~n185 & ~n622;
  assign n624 = ~n126 & n623;
  assign n625 = n524 & n624;
  assign n627 = n61 & n626;
  assign n629 = ~n172 & ~n219;
  assign n630 = ~n628 & n629;
  assign n631 = ~n627 & ~n630;
  assign n632 = n625 & ~n631;
  assign n200 = ~n198 & ~n199;
  assign n633 = n200 & n433;
  assign n634 = ~n173 & ~n186;
  assign n635 = n475 & n634;
  assign n636 = n633 & n635;
  assign n637 = n632 & n636;
  assign n275 = n95 & ~n270;
  assign n641 = n108 & ~n275;
  assign n206 = ~n204 & ~n205;
  assign n643 = ~n174 & n206;
  assign n644 = n642 & n643;
  assign n645 = n641 & n644;
  assign n646 = ~n640 & n645;
  assign n648 = ~n142 & ~n647;
  assign n649 = n526 & n648;
  assign n210 = ~n208 & ~n209;
  assign n242 = n60 & ~n123;
  assign n651 = n210 & ~n242;
  assign n652 = n650 & n651;
  assign n653 = n649 & n652;
  assign n656 = n184 & ~n655;
  assign n657 = ~n93 & ~n656;
  assign n658 = ~n654 & n657;
  assign n660 = ~n460 & ~n465;
  assign n661 = ~n659 & n660;
  assign n662 = n658 & n661;
  assign n663 = n653 & n662;
  assign n664 = n646 & n663;
  assign n665 = n637 & n664;
  assign n666 = n366 & n665;
  assign n767 = n736 ^ n666;
  assign n768 = n666 ^ n532;
  assign n769 = n666 ^ n565;
  assign n770 = n768 & n769;
  assign n771 = n770 ^ n666;
  assign n772 = ~n767 & ~n771;
  assign n773 = n772 ^ n532;
  assign n774 = n773 ^ n765;
  assign n775 = n766 & ~n774;
  assign n776 = n775 ^ n764;
  assign n777 = n776 ^ n753;
  assign n778 = ~n760 & n777;
  assign n779 = n778 ^ n776;
  assign n617 = ~x22 & ~n38;
  assign n618 = n617 ^ x10;
  assign n621 = n620 ^ n618;
  assign n737 = ~n666 & ~n736;
  assign n738 = ~n532 & ~n737;
  assign n739 = n738 ^ n618;
  assign n740 = n621 & n739;
  assign n741 = n740 ^ n620;
  assign n742 = n741 ^ n595;
  assign n743 = ~n318 & n742;
  assign n616 = n590 ^ n570;
  assign n744 = n743 ^ n616;
  assign n780 = n779 ^ n744;
  assign n781 = n595 & ~n616;
  assign n782 = n780 & n781;
  assign n783 = n741 & ~n779;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~n318 & ~n784;
  assign n786 = n779 ^ n741;
  assign n787 = n742 & ~n786;
  assign n788 = ~n318 & n787;
  assign n789 = n788 ^ n779;
  assign n790 = n616 & ~n789;
  assign n791 = ~n785 & ~n790;
  assign n802 = n801 ^ n791;
  assign n813 = ~x22 & ~n34;
  assign n814 = x6 & ~x22;
  assign n815 = ~n813 & ~n814;
  assign n816 = n815 ^ x7;
  assign n985 = ~n318 & ~n816;
  assign n954 = n666 & n736;
  assign n955 = ~n532 & n954;
  assign n956 = n532 & n737;
  assign n957 = ~n955 & ~n956;
  assign n981 = n579 ^ n532;
  assign n982 = ~n957 & ~n981;
  assign n958 = n572 ^ n532;
  assign n983 = n767 & n958;
  assign n984 = ~n982 & ~n983;
  assign n986 = n985 ^ n984;
  assign n894 = ~n363 & ~n622;
  assign n895 = ~n398 & ~n709;
  assign n896 = n894 & n895;
  assign n897 = ~n241 & ~n436;
  assign n898 = ~n525 & ~n654;
  assign n899 = n897 & n898;
  assign n900 = ~n93 & ~n185;
  assign n901 = n315 & n900;
  assign n902 = n899 & n901;
  assign n903 = n896 & n902;
  assign n907 = ~n452 & n906;
  assign n908 = ~n397 & n907;
  assign n841 = ~n554 & ~n676;
  assign n842 = ~n180 & n841;
  assign n843 = ~n198 & n842;
  assign n909 = ~n264 & ~n720;
  assign n910 = n843 & n909;
  assign n911 = n908 & n910;
  assign n912 = n903 & n911;
  assign n913 = ~n125 & ~n416;
  assign n914 = ~n179 & ~n208;
  assign n915 = ~n426 & n914;
  assign n916 = n913 & n915;
  assign n917 = n354 & n916;
  assign n918 = ~n45 & ~n109;
  assign n919 = ~n115 & n918;
  assign n920 = ~n214 & ~n919;
  assign n921 = ~n375 & n920;
  assign n922 = n917 & n921;
  assign n923 = n184 & ~n512;
  assign n924 = ~n628 & ~n923;
  assign n925 = ~n274 & ~n445;
  assign n926 = n924 & n925;
  assign n927 = ~n371 & ~n845;
  assign n928 = ~n126 & ~n174;
  assign n929 = n927 & n928;
  assign n930 = n926 & n929;
  assign n931 = n56 & ~n304;
  assign n932 = ~n92 & n172;
  assign n933 = ~n931 & ~n932;
  assign n934 = n136 ^ n106;
  assign n935 = n551 ^ n60;
  assign n936 = n136 ^ n60;
  assign n937 = n936 ^ n60;
  assign n938 = n935 & n937;
  assign n939 = n938 ^ n60;
  assign n940 = ~n934 & n939;
  assign n941 = n940 ^ n106;
  assign n942 = n933 & ~n941;
  assign n943 = n684 & n942;
  assign n944 = n930 & n943;
  assign n945 = n922 & n944;
  assign n946 = n912 & n945;
  assign n844 = n509 & n843;
  assign n846 = n172 & ~n655;
  assign n847 = ~n207 & ~n846;
  assign n848 = ~n105 & n847;
  assign n849 = ~n845 & n848;
  assign n850 = n101 & ~n172;
  assign n851 = n81 & n166;
  assign n852 = ~n59 & n851;
  assign n853 = ~n850 & ~n852;
  assign n854 = ~n362 & ~n853;
  assign n855 = n136 & n178;
  assign n856 = n95 & ~n855;
  assign n857 = n854 & ~n856;
  assign n858 = n849 & n857;
  assign n859 = n844 & n858;
  assign n860 = ~n840 & n859;
  assign n861 = ~n837 & n860;
  assign n862 = ~n209 & ~n539;
  assign n863 = ~n491 & n862;
  assign n864 = n413 & n863;
  assign n865 = ~n183 & ~n473;
  assign n866 = ~n327 & n865;
  assign n867 = ~n199 & ~n367;
  assign n868 = ~n260 & ~n473;
  assign n869 = n867 & n868;
  assign n870 = n866 & n869;
  assign n871 = n864 & n870;
  assign n225 = ~n86 & ~n106;
  assign n226 = ~n178 & ~n225;
  assign n228 = n109 & ~n141;
  assign n229 = n45 & n228;
  assign n230 = ~n227 & ~n229;
  assign n231 = ~n226 & n230;
  assign n236 = n101 & n136;
  assign n237 = n56 & ~n236;
  assign n238 = ~n235 & ~n237;
  assign n239 = n234 & n238;
  assign n240 = n231 & n239;
  assign n873 = ~n326 & ~n397;
  assign n874 = n872 & n873;
  assign n875 = n480 & n874;
  assign n876 = n240 & n875;
  assign n877 = n871 & n876;
  assign n878 = ~n60 & ~n510;
  assign n879 = ~n347 & ~n878;
  assign n880 = n315 & ~n879;
  assign n881 = n172 & ~n334;
  assign n882 = ~n102 & ~n881;
  assign n271 = n56 & ~n270;
  assign n883 = ~n271 & ~n465;
  assign n884 = n882 & n883;
  assign n885 = n880 & n884;
  assign n243 = n95 & ~n163;
  assign n244 = ~n242 & ~n243;
  assign n886 = n244 & ~n275;
  assign n888 = ~n363 & ~n721;
  assign n889 = ~n887 & n888;
  assign n890 = n886 & n889;
  assign n891 = n885 & n890;
  assign n892 = n877 & n891;
  assign n893 = n861 & n892;
  assign n987 = n946 ^ n893;
  assign n988 = n946 ^ n736;
  assign n989 = n946 ^ n565;
  assign n990 = n988 & n989;
  assign n991 = n990 ^ n946;
  assign n992 = ~n987 & ~n991;
  assign n993 = n992 ^ n736;
  assign n994 = n993 ^ n984;
  assign n995 = n986 & ~n994;
  assign n996 = n995 ^ n985;
  assign n811 = ~x22 & ~n36;
  assign n812 = n811 ^ x8;
  assign n817 = n816 ^ n812;
  assign n979 = ~n318 & ~n817;
  assign n947 = ~n893 & ~n946;
  assign n948 = ~n736 & ~n947;
  assign n980 = n979 ^ n948;
  assign n997 = n996 ^ n980;
  assign n1104 = ~n318 & ~n812;
  assign n1105 = n571 & ~n1104;
  assign n1106 = n812 ^ n318;
  assign n1107 = n1106 ^ n812;
  assign n1108 = n812 ^ n620;
  assign n1109 = n1108 ^ n812;
  assign n1110 = n1107 & ~n1109;
  assign n1111 = n1110 ^ n812;
  assign n1112 = n546 & ~n1111;
  assign n1113 = n1112 ^ n812;
  assign n1114 = ~n1105 & n1113;
  assign n998 = ~n55 & ~n323;
  assign n999 = n81 & n159;
  assign n1000 = ~n368 & ~n999;
  assign n1001 = n115 & ~n1000;
  assign n1002 = ~n998 & ~n1001;
  assign n1003 = ~n721 & ~n1002;
  assign n1004 = n59 & ~n337;
  assign n1005 = ~n56 & ~n1004;
  assign n1006 = ~n141 & ~n1005;
  assign n1007 = ~n260 & ~n554;
  assign n1008 = ~n712 & n1007;
  assign n1009 = ~n360 & n1008;
  assign n1010 = ~n521 & n1009;
  assign n1011 = ~n1006 & n1010;
  assign n1013 = ~n185 & ~n203;
  assign n1014 = ~n1012 & n1013;
  assign n1015 = ~n681 & n1014;
  assign n1016 = n505 & n1015;
  assign n1017 = n874 & n1016;
  assign n1018 = n1011 & n1017;
  assign n1019 = n1003 & n1018;
  assign n1023 = n463 & n1022;
  assign n1024 = n896 & n1023;
  assign n1025 = ~n474 & ~n510;
  assign n1026 = n92 & n136;
  assign n1027 = n86 & ~n1026;
  assign n1028 = n1025 & ~n1027;
  assign n1029 = ~n264 & ~n403;
  assign n1030 = n927 & n1029;
  assign n1031 = n1028 & n1030;
  assign n1032 = n1024 & n1031;
  assign n211 = n59 & ~n159;
  assign n212 = n210 & ~n211;
  assign n213 = n206 & n212;
  assign n215 = ~n101 & n106;
  assign n216 = ~n214 & ~n215;
  assign n221 = ~n219 & ~n220;
  assign n222 = n53 & ~n221;
  assign n223 = n216 & ~n222;
  assign n224 = n213 & n223;
  assign n1033 = ~n355 & ~n711;
  assign n1034 = n306 & n1026;
  assign n1035 = n60 & ~n1034;
  assign n1036 = ~n374 & ~n1035;
  assign n1037 = n1033 & n1036;
  assign n1038 = n244 & n1037;
  assign n1039 = n224 & n1038;
  assign n1040 = n1032 & n1039;
  assign n1041 = n1019 & n1040;
  assign n1042 = n400 & n882;
  assign n1043 = n184 & ~n289;
  assign n1044 = ~n111 & ~n1043;
  assign n1045 = n1042 & n1044;
  assign n1046 = ~n227 & ~n460;
  assign n1047 = n234 & n1046;
  assign n1048 = ~n278 & ~n628;
  assign n1050 = ~n379 & ~n1049;
  assign n1051 = n1048 & n1050;
  assign n1052 = n1047 & n1051;
  assign n1053 = n1045 & n1052;
  assign n1056 = ~n204 & ~n242;
  assign n1057 = n120 & n904;
  assign n1058 = n172 & ~n1057;
  assign n1059 = n1056 & ~n1058;
  assign n1060 = n1055 & n1059;
  assign n1061 = n1053 & n1060;
  assign n1062 = n1003 & n1061;
  assign n1065 = n86 & ~n124;
  assign n1066 = n1064 & ~n1065;
  assign n1067 = n415 & n1066;
  assign n1068 = n865 & n1067;
  assign n1069 = n167 & n346;
  assign n1070 = ~n60 & n1069;
  assign n1071 = n346 & n351;
  assign n1072 = n45 & ~n53;
  assign n1073 = ~n1071 & n1072;
  assign n1074 = ~n1070 & n1073;
  assign n1075 = n95 & ~n335;
  assign n1076 = ~n397 & ~n1075;
  assign n1077 = n101 & n289;
  assign n1078 = n59 & ~n1077;
  assign n1079 = n1076 & ~n1078;
  assign n1080 = n928 & n1079;
  assign n1081 = ~n1074 & n1080;
  assign n1082 = n1068 & n1081;
  assign n1084 = n290 & n1083;
  assign n1085 = ~n55 & ~n95;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = n1082 & ~n1086;
  assign n161 = ~n142 & ~n160;
  assign n168 = n56 & ~n167;
  assign n169 = n161 & ~n168;
  assign n170 = n138 & n169;
  assign n1088 = n110 & ~n1071;
  assign n1089 = ~n443 & ~n1088;
  assign n1090 = n270 & n838;
  assign n1091 = n56 & ~n1090;
  assign n1092 = ~n125 & ~n1091;
  assign n1093 = n1089 & n1092;
  assign n1094 = n170 & n1093;
  assign n1095 = n1087 & n1094;
  assign n1096 = n1062 & n1095;
  assign n1097 = ~n893 & n1096;
  assign n1098 = ~n1041 & n1097;
  assign n1099 = n893 & n1041;
  assign n1100 = n813 ^ x6;
  assign n1101 = ~n318 & n1100;
  assign n1102 = ~n1099 & ~n1101;
  assign n1103 = ~n1098 & ~n1102;
  assign n1115 = n1114 ^ n1103;
  assign n1116 = n618 ^ n558;
  assign n1117 = ~n748 & ~n1116;
  assign n969 = n595 ^ n558;
  assign n1118 = n533 & ~n969;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = n1119 ^ n1103;
  assign n1121 = ~n1115 & ~n1120;
  assign n1122 = n1121 ^ n1119;
  assign n1123 = n1122 ^ n996;
  assign n1124 = ~n997 & n1123;
  assign n1125 = n1124 ^ n1122;
  assign n977 = n773 ^ n766;
  assign n963 = n546 & n621;
  assign n964 = n963 ^ n620;
  assign n965 = ~n571 & n964;
  assign n966 = ~n318 & ~n620;
  assign n967 = ~n965 & ~n966;
  assign n959 = ~n957 & n958;
  assign n960 = n565 ^ n532;
  assign n961 = n767 & n960;
  assign n962 = ~n959 & ~n961;
  assign n968 = n967 ^ n962;
  assign n970 = ~n748 & ~n969;
  assign n971 = n533 & ~n761;
  assign n972 = ~n970 & ~n971;
  assign n973 = n972 ^ n962;
  assign n974 = ~n968 & n973;
  assign n975 = n974 ^ n972;
  assign n949 = n948 ^ n816;
  assign n950 = ~n817 & n949;
  assign n951 = n950 ^ n816;
  assign n952 = ~n318 & ~n951;
  assign n803 = n318 & n571;
  assign n804 = n318 & n546;
  assign n805 = ~n595 & n804;
  assign n806 = ~n803 & ~n805;
  assign n807 = n571 ^ n546;
  assign n808 = n618 & ~n807;
  assign n809 = n808 ^ n546;
  assign n810 = n806 & n809;
  assign n953 = n952 ^ n810;
  assign n976 = n975 ^ n953;
  assign n978 = n977 ^ n976;
  assign n1126 = n1125 ^ n978;
  assign n1127 = n1122 ^ n997;
  assign n1165 = n816 ^ n318;
  assign n1166 = n1165 ^ n546;
  assign n1167 = n1166 ^ n816;
  assign n1168 = n817 ^ n816;
  assign n1169 = n816 ^ n546;
  assign n1170 = n1169 ^ n816;
  assign n1171 = ~n1168 & n1170;
  assign n1172 = n1171 ^ n816;
  assign n1173 = ~n1167 & n1172;
  assign n1174 = n1173 ^ n1165;
  assign n1175 = ~n803 & n1174;
  assign n1156 = n736 & n947;
  assign n1157 = n893 & n946;
  assign n1158 = ~n736 & n1157;
  assign n1159 = ~n1156 & ~n1158;
  assign n1160 = n736 ^ n572;
  assign n1161 = ~n1159 & n1160;
  assign n1162 = n736 ^ n565;
  assign n1163 = n987 & n1162;
  assign n1164 = ~n1161 & ~n1163;
  assign n1176 = n1175 ^ n1164;
  assign n1177 = n620 ^ n558;
  assign n1178 = ~n748 & ~n1177;
  assign n1179 = n533 & ~n1116;
  assign n1180 = ~n1178 & ~n1179;
  assign n1181 = n1180 ^ n1164;
  assign n1182 = n1176 & n1181;
  assign n1183 = n1182 ^ n1180;
  assign n1153 = n993 ^ n985;
  assign n1154 = n1153 ^ n984;
  assign n1152 = n1119 ^ n1115;
  assign n1155 = n1154 ^ n1152;
  assign n1184 = n1183 ^ n1155;
  assign n1128 = ~n1098 & ~n1099;
  assign n1129 = ~n1041 & ~n1096;
  assign n1130 = n893 & n1129;
  assign n1131 = n1041 & n1096;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = ~n565 & ~n1132;
  assign n1134 = n1128 & ~n1133;
  assign n1135 = n1041 & ~n1134;
  assign n29 = ~x22 & ~n28;
  assign n30 = n29 ^ x5;
  assign n1136 = n30 & ~n318;
  assign n1137 = ~n1133 & ~n1136;
  assign n1138 = ~n1135 & ~n1137;
  assign n1139 = ~n1098 & n1138;
  assign n1140 = ~n1101 & n1139;
  assign n1141 = n595 ^ n532;
  assign n1142 = ~n957 & ~n1141;
  assign n1143 = n767 & ~n981;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = n1101 ^ n1099;
  assign n1146 = ~n1138 & n1145;
  assign n1147 = ~n1144 & ~n1146;
  assign n1148 = ~n1140 & ~n1147;
  assign n1149 = ~n1101 & n1144;
  assign n1150 = n1098 & ~n1149;
  assign n1151 = n1148 & ~n1150;
  assign n1185 = n1184 ^ n1151;
  assign n1191 = n736 ^ n579;
  assign n1192 = ~n1159 & ~n1191;
  assign n1193 = n987 & n1160;
  assign n1194 = ~n1192 & ~n1193;
  assign n1187 = n618 ^ n532;
  assign n1188 = ~n957 & ~n1187;
  assign n1189 = n767 & ~n1141;
  assign n1190 = ~n1188 & ~n1189;
  assign n1195 = n1194 ^ n1190;
  assign n1196 = n812 ^ n558;
  assign n1197 = ~n748 & ~n1196;
  assign n1198 = n533 & ~n1177;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = n1199 ^ n1190;
  assign n1201 = ~n1195 & n1200;
  assign n1202 = n1201 ^ n1199;
  assign n1186 = n1180 ^ n1176;
  assign n1203 = n1202 ^ n1186;
  assign n1212 = n736 ^ n595;
  assign n1213 = ~n1159 & ~n1212;
  assign n1214 = n987 & ~n1191;
  assign n1215 = ~n1213 & ~n1214;
  assign n1208 = n620 ^ n532;
  assign n1209 = ~n957 & ~n1208;
  assign n1210 = n767 & ~n1187;
  assign n1211 = ~n1209 & ~n1210;
  assign n1216 = n1215 ^ n1211;
  assign n1217 = n816 ^ n558;
  assign n1218 = ~n748 & n1217;
  assign n1219 = n533 & ~n1196;
  assign n1220 = ~n1218 & ~n1219;
  assign n1221 = n1220 ^ n1211;
  assign n1222 = ~n1216 & n1221;
  assign n1223 = n1222 ^ n1220;
  assign n1204 = n754 & ~n816;
  assign n1205 = n756 & n1100;
  assign n1206 = n1205 ^ n318;
  assign n1207 = ~n1204 & n1206;
  assign n1224 = n1223 ^ n1207;
  assign n31 = ~x22 & ~n27;
  assign n32 = n31 ^ x4;
  assign n1236 = n32 & ~n318;
  assign n1225 = ~n572 & ~n1132;
  assign n1226 = n1041 ^ n893;
  assign n1227 = n1226 ^ n565;
  assign n1228 = n1227 ^ n1096;
  assign n1229 = n1228 ^ n893;
  assign n1230 = n1229 ^ n565;
  assign n1231 = n1097 ^ n893;
  assign n1232 = n1231 ^ n565;
  assign n1233 = ~n1230 & n1232;
  assign n1234 = n1233 ^ n1227;
  assign n1235 = ~n1225 & ~n1234;
  assign n1237 = n1236 ^ n1235;
  assign n1238 = n1236 ^ n1041;
  assign n1239 = ~n1096 & ~n1238;
  assign n1240 = n1239 ^ n1041;
  assign n1241 = ~n1237 & ~n1240;
  assign n1242 = ~n572 & n1130;
  assign n1243 = ~n1236 & ~n1242;
  assign n1244 = n572 & n1097;
  assign n1245 = n1041 & ~n1244;
  assign n1246 = ~n1243 & ~n1245;
  assign n1247 = ~n1241 & ~n1246;
  assign n1248 = n1247 ^ n1207;
  assign n1249 = n1224 & ~n1248;
  assign n1250 = n1249 ^ n1223;
  assign n1251 = n1250 ^ n1202;
  assign n1252 = n1203 & n1251;
  assign n1253 = n1252 ^ n1250;
  assign n1254 = n1253 ^ n1151;
  assign n1255 = ~n1185 & n1254;
  assign n1256 = n1255 ^ n1253;
  assign n1257 = ~n1127 & ~n1256;
  assign n1258 = n1126 & ~n1257;
  assign n1259 = n1250 ^ n1203;
  assign n1260 = ~n893 & n1131;
  assign n1261 = ~n1130 & ~n1260;
  assign n1262 = n893 ^ n30;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n1096 ^ n1041;
  assign n1265 = n1100 ^ n893;
  assign n1266 = n1264 & ~n1265;
  assign n1267 = ~n1263 & ~n1266;
  assign n1281 = ~n275 & n1280;
  assign n1282 = ~n233 & n1056;
  assign n1285 = n1283 & n1284;
  assign n1286 = n1282 & n1285;
  assign n1287 = n490 & n1286;
  assign n1288 = n184 & ~n638;
  assign n1289 = ~n416 & ~n1288;
  assign n1290 = ~n362 & n1289;
  assign n1291 = n163 ^ n60;
  assign n1292 = n163 ^ n136;
  assign n1293 = n1292 ^ n136;
  assign n1294 = n1085 ^ n136;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = n1295 ^ n136;
  assign n1297 = ~n1291 & n1296;
  assign n1298 = n1297 ^ n60;
  assign n1299 = n1290 & ~n1298;
  assign n1300 = n1287 & n1299;
  assign n1301 = n71 & ~n219;
  assign n1302 = ~n45 & ~n1301;
  assign n1303 = ~n94 & ~n1302;
  assign n1304 = ~n918 & ~n1301;
  assign n1305 = n159 & ~n1304;
  assign n1306 = ~n1303 & ~n1305;
  assign n1307 = n106 & ~n427;
  assign n1308 = ~n186 & ~n1307;
  assign n1309 = ~n1306 & n1308;
  assign n1310 = n293 & n1309;
  assign n1311 = n1300 & n1310;
  assign n1312 = n1281 & n1311;
  assign n1313 = n1041 ^ n812;
  assign n1314 = n1313 ^ n816;
  assign n1315 = n1314 ^ n1313;
  assign n1316 = n1313 ^ n812;
  assign n1317 = n1315 & ~n1316;
  assign n1318 = n1317 ^ n1313;
  assign n1319 = n1312 & ~n1318;
  assign n1320 = n1319 ^ n1313;
  assign n1321 = ~n1267 & ~n1320;
  assign n1322 = ~x22 & ~n26;
  assign n1323 = n1322 ^ x3;
  assign n1324 = n987 & n1323;
  assign n1325 = n948 & ~n1324;
  assign n1326 = n736 ^ n32;
  assign n1327 = n987 & ~n1326;
  assign n1328 = n1323 ^ n1156;
  assign n1329 = n1328 ^ n1156;
  assign n1330 = n1158 ^ n1156;
  assign n1331 = ~n1329 & n1330;
  assign n1332 = n1331 ^ n1156;
  assign n1333 = ~n1327 & ~n1332;
  assign n1334 = n1325 & ~n1333;
  assign n1335 = n1321 & n1334;
  assign n1336 = n767 & n1323;
  assign n1337 = n1320 ^ n1267;
  assign n1338 = ~n1325 & n1333;
  assign n1339 = n1338 ^ n1320;
  assign n1340 = n1337 & ~n1339;
  assign n1341 = n1340 ^ n1267;
  assign n1342 = n1336 & ~n1341;
  assign n1343 = ~n1335 & ~n1342;
  assign n1348 = ~n1159 & ~n1326;
  assign n1349 = n736 ^ n30;
  assign n1350 = n987 & ~n1349;
  assign n1351 = ~n1348 & ~n1350;
  assign n1344 = ~n1261 & ~n1265;
  assign n1345 = n893 ^ n816;
  assign n1346 = n1264 & n1345;
  assign n1347 = ~n1344 & ~n1346;
  assign n1352 = n1351 ^ n1347;
  assign n1353 = n1041 ^ n620;
  assign n1354 = n1353 ^ n812;
  assign n1355 = n1354 ^ n1353;
  assign n1356 = n1353 ^ n620;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = n1357 ^ n1353;
  assign n1359 = n1312 & ~n1358;
  assign n1360 = n1359 ^ n1353;
  assign n1361 = n1360 ^ n1351;
  assign n1362 = n1352 & ~n1361;
  assign n1363 = n1362 ^ n1347;
  assign n1364 = n1343 & n1363;
  assign n1408 = ~n1261 & n1345;
  assign n1365 = n893 ^ n812;
  assign n1409 = n1264 & ~n1365;
  assign n1410 = ~n1408 & ~n1409;
  assign n1405 = ~n1159 & ~n1349;
  assign n1379 = n1100 ^ n736;
  assign n1406 = n987 & ~n1379;
  assign n1407 = ~n1405 & ~n1406;
  assign n1411 = n1410 ^ n1407;
  assign n1397 = n532 ^ n32;
  assign n1412 = n767 & ~n1397;
  assign n1413 = n956 ^ n955;
  assign n1414 = n1323 ^ n955;
  assign n1415 = n1414 ^ n955;
  assign n1416 = n1413 & n1415;
  assign n1417 = n1416 ^ n955;
  assign n1418 = ~n1412 & ~n1417;
  assign n1419 = n1418 ^ n1410;
  assign n1420 = n1411 & ~n1419;
  assign n1421 = n1420 ^ n1407;
  assign n1402 = n533 & n1323;
  assign n1398 = ~n957 & ~n1397;
  assign n1399 = n532 ^ n30;
  assign n1400 = n767 & ~n1399;
  assign n1401 = ~n1398 & ~n1400;
  assign n1403 = n1402 ^ n1401;
  assign n1385 = n738 & ~n1323;
  assign n1386 = ~n955 & ~n1385;
  assign n1387 = n1041 ^ n618;
  assign n1388 = n1387 ^ n620;
  assign n1389 = n1388 ^ n1387;
  assign n1390 = n1387 ^ n618;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = n1391 ^ n1387;
  assign n1393 = n1312 & ~n1392;
  assign n1394 = n1393 ^ n1387;
  assign n1395 = ~n1386 & ~n1394;
  assign n1380 = ~n1159 & ~n1379;
  assign n1381 = n816 ^ n736;
  assign n1382 = n987 & n1381;
  assign n1383 = ~n1380 & ~n1382;
  assign n1370 = n1041 ^ n595;
  assign n1371 = n1370 ^ n618;
  assign n1372 = n1371 ^ n1370;
  assign n1373 = n1370 ^ n595;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = n1374 ^ n1370;
  assign n1376 = n1312 & ~n1375;
  assign n1377 = n1376 ^ n1370;
  assign n1366 = ~n1261 & ~n1365;
  assign n1367 = n893 ^ n620;
  assign n1368 = n1264 & ~n1367;
  assign n1369 = ~n1366 & ~n1368;
  assign n1378 = n1377 ^ n1369;
  assign n1384 = n1383 ^ n1378;
  assign n1396 = n1395 ^ n1384;
  assign n1404 = n1403 ^ n1396;
  assign n1422 = n1421 ^ n1404;
  assign n1423 = ~n1364 & ~n1422;
  assign n1425 = n1341 ^ n1336;
  assign n1426 = n1425 ^ n1321;
  assign n1427 = ~n1334 & n1426;
  assign n1428 = n1427 ^ n1321;
  assign n1424 = n1360 ^ n1352;
  assign n1429 = n1428 ^ n1424;
  assign n1434 = n1041 ^ n816;
  assign n1435 = n1434 ^ n1100;
  assign n1436 = n1435 ^ n1434;
  assign n1437 = n1434 ^ n816;
  assign n1438 = ~n1436 & ~n1437;
  assign n1439 = n1438 ^ n1434;
  assign n1440 = n1312 & n1439;
  assign n1441 = n1440 ^ n1434;
  assign n1430 = n893 ^ n32;
  assign n1431 = ~n1261 & ~n1430;
  assign n1432 = ~n1262 & n1264;
  assign n1433 = ~n1431 & ~n1432;
  assign n1442 = n1441 ^ n1433;
  assign n1443 = n1323 ^ n1096;
  assign n1444 = n1264 & ~n1443;
  assign n1445 = n1444 ^ n1096;
  assign n1446 = ~n893 & n1445;
  assign n1447 = ~n1324 & ~n1446;
  assign n1448 = ~n1442 & ~n1447;
  assign n1449 = n1100 ^ n1041;
  assign n1450 = n1449 ^ n1100;
  assign n1451 = n1100 ^ n30;
  assign n1452 = n1451 ^ n1100;
  assign n1453 = ~n1450 & n1452;
  assign n1454 = n1453 ^ n1100;
  assign n1455 = n1312 & n1454;
  assign n1456 = n1455 ^ n1449;
  assign n1457 = ~n1448 & n1456;
  assign n1458 = n1264 & ~n1430;
  assign n1459 = n1260 ^ n1130;
  assign n1460 = n1323 ^ n1260;
  assign n1461 = n1460 ^ n1260;
  assign n1462 = n1459 & n1461;
  assign n1463 = n1462 ^ n1260;
  assign n1464 = ~n1458 & ~n1463;
  assign n1465 = n1442 & n1464;
  assign n1466 = ~n1446 & n1465;
  assign n1467 = ~n1457 & ~n1466;
  assign n1468 = ~n1442 & ~n1464;
  assign n1469 = ~n1324 & ~n1468;
  assign n1470 = n1467 & ~n1469;
  assign n1472 = n30 & ~n1312;
  assign n1471 = ~n1096 & n1323;
  assign n1473 = n1472 ^ n1471;
  assign n1474 = n1323 ^ n1312;
  assign n1475 = n1312 ^ n1041;
  assign n1476 = ~n1312 & n1475;
  assign n1477 = n1476 ^ n1312;
  assign n1478 = ~n1474 & ~n1477;
  assign n1479 = n1478 ^ n1476;
  assign n1480 = n1479 ^ n1312;
  assign n1481 = n1480 ^ n1041;
  assign n1482 = n32 & n1481;
  assign n1483 = n1482 ^ n1041;
  assign n1484 = n1483 ^ n1472;
  assign n1485 = n1484 ^ n1483;
  assign n1486 = n1483 ^ n1041;
  assign n1487 = n1485 & ~n1486;
  assign n1488 = n1487 ^ n1483;
  assign n1489 = ~n1473 & ~n1488;
  assign n1490 = ~n1470 & ~n1489;
  assign n1491 = ~n1465 & ~n1469;
  assign n1492 = n1456 & ~n1491;
  assign n1493 = n1333 ^ n1325;
  assign n1494 = n1493 ^ n1337;
  assign n1495 = n1494 ^ n1447;
  assign n1496 = n1494 ^ n1441;
  assign n1497 = n1494 ^ n1442;
  assign n1498 = n1494 & n1497;
  assign n1499 = n1498 ^ n1494;
  assign n1500 = ~n1496 & n1499;
  assign n1501 = n1500 ^ n1498;
  assign n1502 = n1501 ^ n1494;
  assign n1503 = n1502 ^ n1442;
  assign n1504 = n1495 & n1503;
  assign n1505 = n1504 ^ n1494;
  assign n1506 = ~n1492 & ~n1505;
  assign n1507 = ~n1490 & n1506;
  assign n1508 = n1507 ^ n1424;
  assign n1509 = n1508 ^ n1424;
  assign n1510 = n1446 & ~n1456;
  assign n1511 = n1510 ^ n1441;
  assign n1512 = ~n1442 & ~n1511;
  assign n1513 = n1512 ^ n1433;
  assign n1514 = ~n1494 & ~n1513;
  assign n1515 = n1514 ^ n1424;
  assign n1516 = n1515 ^ n1424;
  assign n1517 = ~n1509 & ~n1516;
  assign n1518 = n1517 ^ n1424;
  assign n1519 = n1429 & ~n1518;
  assign n1520 = n1519 ^ n1428;
  assign n1521 = ~n1423 & n1520;
  assign n1522 = ~n1343 & ~n1363;
  assign n1523 = n1422 & ~n1522;
  assign n1524 = n1394 ^ n1386;
  assign n1525 = n1418 ^ n1411;
  assign n1526 = ~n1524 & n1525;
  assign n1527 = ~n1523 & ~n1526;
  assign n1528 = ~n1521 & n1527;
  assign n1529 = n1524 & ~n1525;
  assign n1530 = n1529 ^ n1422;
  assign n1531 = n1363 ^ n1343;
  assign n1532 = n1520 ^ n1363;
  assign n1533 = n1531 & ~n1532;
  assign n1534 = n1533 ^ n1343;
  assign n1535 = n1534 ^ n1529;
  assign n1536 = ~n1530 & n1535;
  assign n1537 = n1536 ^ n1422;
  assign n1538 = ~n1528 & n1537;
  assign n1547 = ~n1261 & ~n1367;
  assign n1548 = n893 ^ n618;
  assign n1549 = n1264 & ~n1548;
  assign n1550 = ~n1547 & ~n1549;
  assign n1543 = ~n1159 & n1381;
  assign n1544 = n812 ^ n736;
  assign n1545 = n987 & ~n1544;
  assign n1546 = ~n1543 & ~n1545;
  assign n1551 = n1550 ^ n1546;
  assign n1539 = ~n957 & ~n1399;
  assign n1540 = n1100 ^ n532;
  assign n1541 = n767 & ~n1540;
  assign n1542 = ~n1539 & ~n1541;
  assign n1552 = n1551 ^ n1542;
  assign n1553 = n1538 & n1552;
  assign n1612 = n1546 ^ n1542;
  assign n1613 = ~n1551 & n1612;
  assign n1614 = n1613 ^ n1542;
  assign n1610 = n754 & n1323;
  assign n1557 = n1041 ^ n579;
  assign n1558 = n1557 ^ n595;
  assign n1559 = n1558 ^ n1557;
  assign n1560 = n1557 ^ n579;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = n1561 ^ n1557;
  assign n1563 = n1312 & ~n1562;
  assign n1564 = n1563 ^ n1557;
  assign n1565 = n593 & ~n1402;
  assign n1608 = ~n1564 & n1565;
  assign n1603 = ~n1159 & ~n1544;
  assign n1604 = n736 ^ n620;
  assign n1605 = n987 & ~n1604;
  assign n1606 = ~n1603 & ~n1605;
  assign n1599 = ~n957 & ~n1540;
  assign n1600 = n816 ^ n532;
  assign n1601 = n767 & n1600;
  assign n1602 = ~n1599 & ~n1601;
  assign n1607 = n1606 ^ n1602;
  assign n1609 = n1608 ^ n1607;
  assign n1611 = n1610 ^ n1609;
  assign n1615 = n1614 ^ n1611;
  assign n1567 = n558 ^ n32;
  assign n1568 = n533 & ~n1567;
  assign n1569 = n1323 ^ n745;
  assign n1570 = n1569 ^ n745;
  assign n1571 = n747 ^ n745;
  assign n1572 = ~n1570 & n1571;
  assign n1573 = n1572 ^ n745;
  assign n1574 = ~n1568 & ~n1573;
  assign n1566 = n1565 ^ n1564;
  assign n1575 = n1574 ^ n1566;
  assign n1554 = n1383 ^ n1377;
  assign n1555 = n1378 & ~n1554;
  assign n1556 = n1555 ^ n1369;
  assign n1595 = n1574 ^ n1556;
  assign n1596 = ~n1575 & n1595;
  assign n1597 = n1596 ^ n1556;
  assign n1585 = n1041 ^ n572;
  assign n1586 = n1585 ^ n579;
  assign n1587 = n1586 ^ n1585;
  assign n1588 = n1585 ^ n572;
  assign n1589 = ~n1587 & ~n1588;
  assign n1590 = n1589 ^ n1585;
  assign n1591 = n1312 & n1590;
  assign n1592 = n1591 ^ n1585;
  assign n1581 = ~n1261 & ~n1548;
  assign n1582 = n893 ^ n595;
  assign n1583 = n1264 & ~n1582;
  assign n1584 = ~n1581 & ~n1583;
  assign n1593 = n1592 ^ n1584;
  assign n1577 = ~n748 & ~n1567;
  assign n1578 = n558 ^ n30;
  assign n1579 = n533 & ~n1578;
  assign n1580 = ~n1577 & ~n1579;
  assign n1594 = n1593 ^ n1580;
  assign n1598 = n1597 ^ n1594;
  assign n1616 = n1615 ^ n1598;
  assign n1576 = n1575 ^ n1556;
  assign n1617 = n1616 ^ n1576;
  assign n1618 = n1384 & n1421;
  assign n1619 = n1401 ^ n1395;
  assign n1620 = n1403 & ~n1619;
  assign n1621 = n1620 ^ n1395;
  assign n1622 = n1618 & ~n1621;
  assign n1623 = ~n1384 & ~n1421;
  assign n1624 = n1401 & ~n1402;
  assign n1625 = ~n1395 & n1624;
  assign n1626 = ~n1623 & n1625;
  assign n1627 = ~n1622 & ~n1626;
  assign n1628 = n1627 ^ n1616;
  assign n1629 = n1628 ^ n1627;
  assign n1630 = n1621 & n1623;
  assign n1631 = ~n1401 & n1402;
  assign n1632 = n1395 & n1631;
  assign n1633 = ~n1618 & n1632;
  assign n1634 = ~n1630 & ~n1633;
  assign n1635 = n1634 ^ n1627;
  assign n1636 = ~n1629 & n1635;
  assign n1637 = n1636 ^ n1627;
  assign n1638 = ~n1617 & n1637;
  assign n1639 = n1638 ^ n1576;
  assign n1640 = ~n1553 & ~n1639;
  assign n1641 = ~n1576 & n1627;
  assign n1642 = n1634 & ~n1641;
  assign n1643 = n1642 ^ n1616;
  assign n1644 = n1642 ^ n1552;
  assign n1645 = n1644 ^ n1642;
  assign n1646 = n1642 ^ n1538;
  assign n1647 = n1646 ^ n1642;
  assign n1648 = ~n1645 & ~n1647;
  assign n1649 = n1648 ^ n1642;
  assign n1650 = ~n1643 & n1649;
  assign n1651 = n1650 ^ n1616;
  assign n1652 = ~n1640 & ~n1651;
  assign n1666 = n1323 ^ n318;
  assign n1667 = n1666 ^ n546;
  assign n1668 = n1667 ^ n1666;
  assign n1669 = n1666 ^ n32;
  assign n1670 = n1669 ^ n1666;
  assign n1671 = n1668 & n1670;
  assign n1672 = n1671 ^ n1666;
  assign n1673 = ~n756 & ~n1672;
  assign n1674 = n1673 ^ n1666;
  assign n1675 = ~n803 & ~n1674;
  assign n1657 = n1041 ^ n565;
  assign n1658 = n1657 ^ n572;
  assign n1659 = n1658 ^ n1657;
  assign n1660 = n1657 ^ n565;
  assign n1661 = n1659 & ~n1660;
  assign n1662 = n1661 ^ n1657;
  assign n1663 = n1312 & n1662;
  assign n1664 = n1663 ^ n1657;
  assign n1665 = n1664 ^ n318;
  assign n1676 = n1675 ^ n1665;
  assign n1653 = ~n1261 & ~n1582;
  assign n1654 = n893 ^ n579;
  assign n1655 = n1264 & ~n1654;
  assign n1656 = ~n1653 & ~n1655;
  assign n1677 = n1676 ^ n1656;
  assign n1678 = n1615 ^ n1594;
  assign n1679 = ~n1598 & n1678;
  assign n1680 = n1679 ^ n1597;
  assign n1681 = ~n1677 & n1680;
  assign n1735 = n1608 ^ n1606;
  assign n1736 = n1607 & n1735;
  assign n1737 = n1736 ^ n1602;
  assign n1700 = ~n748 & ~n1578;
  assign n1701 = n1100 ^ n558;
  assign n1702 = n533 & ~n1701;
  assign n1703 = ~n1700 & ~n1702;
  assign n1695 = ~n1159 & ~n1604;
  assign n1696 = n736 ^ n618;
  assign n1697 = n987 & ~n1696;
  assign n1698 = ~n1695 & ~n1697;
  assign n1691 = ~n957 & n1600;
  assign n1692 = n812 ^ n532;
  assign n1693 = n767 & ~n1692;
  assign n1694 = ~n1691 & ~n1693;
  assign n1699 = n1698 ^ n1694;
  assign n1734 = n1703 ^ n1699;
  assign n1738 = n1737 ^ n1734;
  assign n1739 = n1584 ^ n1580;
  assign n1740 = n1593 & n1739;
  assign n1741 = n1740 ^ n1580;
  assign n1742 = n1741 ^ n1734;
  assign n1743 = n1738 & ~n1742;
  assign n1744 = n1743 ^ n1737;
  assign n1727 = ~n1159 & ~n1696;
  assign n1728 = n987 & ~n1212;
  assign n1729 = ~n1727 & ~n1728;
  assign n1724 = ~n957 & ~n1692;
  assign n1725 = n767 & ~n1208;
  assign n1726 = ~n1724 & ~n1725;
  assign n1730 = n1729 ^ n1726;
  assign n1721 = ~n748 & ~n1701;
  assign n1722 = n533 & n1217;
  assign n1723 = ~n1721 & ~n1722;
  assign n1731 = n1730 ^ n1723;
  assign n1717 = n1665 ^ n1656;
  assign n1718 = n1676 & n1717;
  assign n1719 = n1718 ^ n1656;
  assign n1713 = ~n565 & n1312;
  assign n1714 = ~n1041 & ~n1713;
  assign n1712 = ~n318 & n1323;
  assign n1715 = n1714 ^ n1712;
  assign n1708 = ~n1261 & ~n1654;
  assign n1709 = n893 ^ n572;
  assign n1710 = n1264 & n1709;
  assign n1711 = ~n1708 & ~n1710;
  assign n1716 = n1715 ^ n1711;
  assign n1720 = n1719 ^ n1716;
  assign n1732 = n1731 ^ n1720;
  assign n1704 = n1703 ^ n1694;
  assign n1705 = ~n1699 & n1704;
  assign n1706 = n1705 ^ n1703;
  assign n1683 = ~n32 & ~n318;
  assign n1684 = n571 & ~n1683;
  assign n1685 = ~n30 & n318;
  assign n1686 = n1685 ^ n32;
  assign n1687 = n546 & ~n1686;
  assign n1688 = n1687 ^ n32;
  assign n1689 = ~n1684 & n1688;
  assign n1682 = ~n318 & n1664;
  assign n1690 = n1689 ^ n1682;
  assign n1707 = n1706 ^ n1690;
  assign n1733 = n1732 ^ n1707;
  assign n1745 = n1744 ^ n1733;
  assign n1746 = ~n1681 & ~n1745;
  assign n1747 = n1652 & ~n1746;
  assign n1748 = n1677 & ~n1680;
  assign n1749 = n1745 & ~n1748;
  assign n1750 = n1741 ^ n1738;
  assign n1751 = n1614 ^ n1610;
  assign n1752 = n1611 & n1751;
  assign n1753 = n1752 ^ n1609;
  assign n1754 = n1750 & ~n1753;
  assign n1755 = ~n1749 & ~n1754;
  assign n1756 = ~n1747 & n1755;
  assign n1757 = ~n1750 & n1753;
  assign n1758 = n1757 ^ n1745;
  assign n1759 = n1680 ^ n1652;
  assign n1760 = n1680 ^ n1677;
  assign n1761 = n1759 & n1760;
  assign n1762 = n1761 ^ n1652;
  assign n1763 = n1762 ^ n1745;
  assign n1764 = ~n1758 & n1763;
  assign n1765 = n1764 ^ n1745;
  assign n1766 = ~n1756 & n1765;
  assign n1767 = n1731 ^ n1716;
  assign n1768 = n1720 & ~n1767;
  assign n1769 = n1768 ^ n1719;
  assign n1770 = ~n1766 & ~n1769;
  assign n1787 = n1220 ^ n1216;
  assign n1788 = n1787 ^ n1237;
  assign n1784 = n1706 ^ n1682;
  assign n1785 = ~n1690 & ~n1784;
  assign n1786 = n1785 ^ n1706;
  assign n1789 = n1788 ^ n1786;
  assign n1778 = n1712 ^ n1711;
  assign n1779 = n1714 ^ n1711;
  assign n1780 = ~n1778 & n1779;
  assign n1781 = n1780 ^ n1712;
  assign n1774 = n754 & n1100;
  assign n1775 = n30 & n756;
  assign n1776 = n1775 ^ n318;
  assign n1777 = ~n1774 & n1776;
  assign n1782 = n1781 ^ n1777;
  assign n1771 = n1726 ^ n1723;
  assign n1772 = ~n1730 & n1771;
  assign n1773 = n1772 ^ n1723;
  assign n1783 = n1782 ^ n1773;
  assign n1790 = n1789 ^ n1783;
  assign n1791 = n1744 ^ n1707;
  assign n1792 = ~n1733 & n1791;
  assign n1793 = n1792 ^ n1744;
  assign n1794 = n1793 ^ n1783;
  assign n1795 = ~n1790 & n1794;
  assign n1805 = n1787 ^ n1786;
  assign n1806 = n1788 & n1805;
  assign n1807 = n1806 ^ n1786;
  assign n1803 = n1247 ^ n1224;
  assign n1799 = n1777 ^ n1773;
  assign n1800 = ~n1782 & ~n1799;
  assign n1801 = n1800 ^ n1781;
  assign n1797 = n1136 ^ n1134;
  assign n1796 = n1199 ^ n1195;
  assign n1798 = n1797 ^ n1796;
  assign n1802 = n1801 ^ n1798;
  assign n1804 = n1803 ^ n1802;
  assign n1808 = n1807 ^ n1804;
  assign n1809 = n1808 ^ n1789;
  assign n1810 = n1795 & ~n1809;
  assign n1811 = n1810 ^ n1808;
  assign n1812 = ~n1770 & n1811;
  assign n1814 = ~n1790 & ~n1794;
  assign n1815 = n1814 ^ n1793;
  assign n1813 = n1766 & n1769;
  assign n1816 = n1815 ^ n1813;
  assign n1817 = n1815 ^ n1808;
  assign n1818 = n1816 & n1817;
  assign n1819 = n1818 ^ n1815;
  assign n1820 = ~n1812 & ~n1819;
  assign n1821 = n1259 & n1820;
  assign n1826 = n1144 ^ n1101;
  assign n1825 = ~n1099 & ~n1139;
  assign n1827 = n1826 ^ n1825;
  assign n1822 = n1801 ^ n1796;
  assign n1823 = n1798 & ~n1822;
  assign n1824 = n1823 ^ n1801;
  assign n1828 = n1827 ^ n1824;
  assign n1829 = n1807 ^ n1802;
  assign n1830 = ~n1804 & n1829;
  assign n1831 = n1830 ^ n1807;
  assign n1832 = n1831 ^ n1827;
  assign n1833 = n1828 & ~n1832;
  assign n1834 = n1253 ^ n1185;
  assign n1835 = n1834 ^ n1824;
  assign n1836 = n1833 & ~n1835;
  assign n1837 = n1836 ^ n1834;
  assign n1838 = ~n1821 & n1837;
  assign n1840 = n1831 ^ n1824;
  assign n1841 = n1828 & ~n1840;
  assign n1842 = n1841 ^ n1831;
  assign n1839 = ~n1259 & ~n1820;
  assign n1843 = n1842 ^ n1839;
  assign n1844 = n1842 ^ n1834;
  assign n1845 = n1843 & n1844;
  assign n1846 = n1845 ^ n1842;
  assign n1847 = ~n1838 & ~n1846;
  assign n1848 = ~n1258 & n1847;
  assign n1849 = n972 ^ n968;
  assign n1850 = n1183 ^ n1154;
  assign n1851 = n1155 & ~n1850;
  assign n1852 = n1851 ^ n1152;
  assign n1853 = ~n1849 & ~n1852;
  assign n1854 = n1127 & n1256;
  assign n1855 = ~n1126 & ~n1854;
  assign n1856 = ~n1853 & ~n1855;
  assign n1857 = ~n1848 & n1856;
  assign n1858 = n1849 & n1852;
  assign n1859 = n1858 ^ n1126;
  assign n1860 = n1256 ^ n1127;
  assign n1861 = n1847 ^ n1256;
  assign n1862 = n1860 & n1861;
  assign n1863 = n1862 ^ n1127;
  assign n1864 = n1863 ^ n1126;
  assign n1865 = n1859 & ~n1864;
  assign n1866 = n1865 ^ n1858;
  assign n1867 = ~n1857 & ~n1866;
  assign n1868 = ~n318 & n621;
  assign n1869 = n1868 ^ n738;
  assign n1870 = n776 ^ n760;
  assign n1871 = n975 ^ n952;
  assign n1872 = ~n953 & ~n1871;
  assign n1873 = n1872 ^ n975;
  assign n1874 = n1870 & n1873;
  assign n1875 = n1869 & n1874;
  assign n1876 = n1125 ^ n976;
  assign n1877 = ~n978 & n1876;
  assign n1878 = n1877 ^ n1125;
  assign n1879 = ~n1875 & ~n1878;
  assign n1880 = n1873 ^ n1870;
  assign n1881 = n1873 ^ n1869;
  assign n1882 = n1880 & ~n1881;
  assign n1883 = n1882 ^ n1870;
  assign n1884 = ~n1879 & n1883;
  assign n1885 = ~n1870 & ~n1873;
  assign n1886 = ~n1869 & n1885;
  assign n1887 = ~n1878 & n1886;
  assign n1888 = n780 & ~n1887;
  assign n1889 = ~n1884 & ~n1888;
  assign n1890 = ~n1867 & ~n1889;
  assign n1891 = n1878 & ~n1886;
  assign n1892 = ~n1883 & ~n1891;
  assign n1893 = n1875 & n1878;
  assign n1894 = ~n780 & ~n1893;
  assign n1895 = ~n1892 & ~n1894;
  assign n1896 = ~n1890 & ~n1895;
  assign n1897 = n1896 ^ n791;
  assign n1898 = ~n802 & ~n1897;
  assign n1899 = n1898 ^ n1896;
  assign n610 = ~n546 & ~n565;
  assign n611 = ~n579 & ~n595;
  assign n612 = n611 ^ n573;
  assign n613 = ~n318 & n612;
  assign n614 = ~n610 & ~n613;
  assign n608 = ~n606 & ~n607;
  assign n609 = ~n603 & n608;
  assign n615 = n614 ^ n609;
  assign n1900 = n1899 ^ n615;
  assign n1940 = n1939 ^ n1900;
  assign n1948 = ~n172 & n667;
  assign n1949 = ~n71 & ~n1948;
  assign n1950 = n1912 & ~n1949;
  assign n1951 = n60 & ~n339;
  assign n1952 = n1934 & ~n1951;
  assign n1953 = n106 & ~n336;
  assign n1954 = n1952 & ~n1953;
  assign n1955 = n104 & n1954;
  assign n1956 = n1950 & n1955;
  assign n1957 = ~n204 & ~n241;
  assign n1958 = n415 & n1957;
  assign n1959 = n888 & n1958;
  assign n1960 = n1956 & n1959;
  assign n1961 = ~n214 & ~n676;
  assign n1962 = ~n232 & n1961;
  assign n1963 = ~n267 & ~n501;
  assign n1964 = n55 & n390;
  assign n1965 = n1963 & ~n1964;
  assign n1966 = ~n197 & ~n229;
  assign n1967 = n1965 & n1966;
  assign n1968 = n1962 & n1967;
  assign n1969 = n184 & ~n424;
  assign n1970 = n406 & ~n1969;
  assign n1971 = n1968 & n1970;
  assign n1972 = n477 & n1971;
  assign n1973 = ~n242 & n466;
  assign n1974 = ~n298 & ~n647;
  assign n1975 = n1973 & n1974;
  assign n1976 = n463 & n1975;
  assign n1983 = ~n384 & n1982;
  assign n1984 = n1976 & n1983;
  assign n1985 = n1972 & n1984;
  assign n1986 = n1960 & n1985;
  assign n1942 = ~n1887 & ~n1893;
  assign n1943 = n1892 ^ n1884;
  assign n1944 = ~n1867 & n1943;
  assign n1945 = n1944 ^ n1892;
  assign n1946 = n1942 & ~n1945;
  assign n1947 = n1946 ^ n780;
  assign n1987 = n1986 ^ n1947;
  assign n1991 = n184 & ~n346;
  assign n1992 = ~n116 & ~n1991;
  assign n1993 = n1960 & n1992;
  assign n1995 = n59 & ~n136;
  assign n1996 = ~n521 & ~n1995;
  assign n1997 = n244 & n1996;
  assign n1998 = n1994 & n1997;
  assign n1999 = ~n397 & ~n687;
  assign n2000 = ~n60 & n1999;
  assign n2001 = ~n309 & ~n2000;
  assign n2002 = ~n709 & ~n2001;
  assign n2003 = n1998 & n2002;
  assign n2004 = ~n45 & ~n708;
  assign n2005 = n515 & ~n2004;
  assign n2006 = ~n55 & ~n374;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = ~n183 & ~n2007;
  assign n2009 = n94 & ~n178;
  assign n2010 = n219 ^ n110;
  assign n2011 = n110 ^ n106;
  assign n2012 = n2011 ^ n106;
  assign n2013 = n1034 ^ n106;
  assign n2014 = n2012 & n2013;
  assign n2015 = n2014 ^ n106;
  assign n2016 = n2010 & ~n2015;
  assign n2017 = n2016 ^ n219;
  assign n2018 = ~n2009 & ~n2017;
  assign n2019 = n2008 & n2018;
  assign n2020 = n1931 & n2019;
  assign n2021 = n2003 & n2020;
  assign n2022 = n1993 & n2021;
  assign n1988 = n1880 ^ n1869;
  assign n1989 = n1988 ^ n1878;
  assign n1990 = n1989 ^ n1867;
  assign n2023 = n2022 ^ n1990;
  assign n2056 = n1127 & n1858;
  assign n2057 = ~n1127 & n1853;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n1860 & ~n2058;
  assign n2060 = ~n1256 & ~n2056;
  assign n2061 = n1852 ^ n1849;
  assign n2062 = n1852 ^ n1127;
  assign n2063 = ~n2061 & n2062;
  assign n2064 = n2063 ^ n1127;
  assign n2065 = ~n2060 & n2064;
  assign n2066 = n2065 ^ n1847;
  assign n2067 = n2066 ^ n2065;
  assign n2068 = ~n1256 & ~n2064;
  assign n2069 = ~n2057 & ~n2068;
  assign n2070 = n2069 ^ n2065;
  assign n2071 = n2067 & ~n2070;
  assign n2072 = n2071 ^ n2065;
  assign n2073 = ~n2059 & ~n2072;
  assign n2074 = n2073 ^ n1126;
  assign n2031 = ~n95 & ~n451;
  assign n2032 = ~n115 & ~n2031;
  assign n2033 = ~n166 & n368;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = ~n242 & n2034;
  assign n2036 = ~n362 & ~n506;
  assign n2037 = ~n525 & n2036;
  assign n2038 = n2035 & n2037;
  assign n2039 = ~n241 & ~n319;
  assign n2040 = ~n443 & n2039;
  assign n2041 = n101 & ~n219;
  assign n2042 = ~n110 & n2041;
  assign n2043 = ~n385 & ~n2042;
  assign n2044 = ~n186 & ~n278;
  assign n2045 = ~n676 & n2044;
  assign n2046 = ~n453 & n2045;
  assign n2047 = ~n2043 & n2046;
  assign n2048 = n2040 & n2047;
  assign n2049 = n2038 & n2048;
  assign n2050 = ~n82 & n1072;
  assign n2051 = ~n398 & ~n2050;
  assign n2052 = ~n107 & n2051;
  assign n2053 = n2049 & n2052;
  assign n2054 = n877 & n2053;
  assign n2055 = n2030 & n2054;
  assign n2075 = n2074 ^ n2055;
  assign n2101 = n2061 ^ n1860;
  assign n2102 = n2101 ^ n1847;
  assign n2089 = ~n667 & ~n2088;
  assign n2090 = n2086 & ~n2089;
  assign n2091 = n843 & n2090;
  assign n2092 = n2084 & n2091;
  assign n2093 = n110 & ~n309;
  assign n2094 = ~n465 & ~n2093;
  assign n2095 = n234 & n2094;
  assign n2096 = n857 & n2095;
  assign n2097 = n907 & n2096;
  assign n2098 = n2092 & n2097;
  assign n2099 = n330 & n903;
  assign n2100 = n2098 & n2099;
  assign n2103 = n2102 ^ n2100;
  assign n130 = ~n92 & ~n129;
  assign n181 = ~n179 & ~n180;
  assign n182 = n175 & n181;
  assign n187 = ~n159 & n184;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~n185 & n188;
  assign n190 = ~n183 & n189;
  assign n191 = n182 & n190;
  assign n192 = n170 & n191;
  assign n193 = ~n130 & n192;
  assign n194 = n104 & n193;
  assign n201 = ~n197 & n200;
  assign n202 = n194 & n201;
  assign n2110 = ~n355 & ~n416;
  assign n2111 = ~n319 & ~n507;
  assign n2112 = n2110 & n2111;
  assign n257 = n71 & n256;
  assign n258 = n86 & ~n257;
  assign n259 = ~n255 & ~n258;
  assign n2113 = n259 & ~n375;
  assign n2114 = n2112 & n2113;
  assign n2115 = ~n209 & ~n453;
  assign n2116 = ~n501 & n2115;
  assign n2117 = n2114 & n2116;
  assign n2118 = n875 & n2117;
  assign n2119 = ~n510 & ~n721;
  assign n2120 = ~n294 & n2119;
  assign n2121 = ~n232 & ~n622;
  assign n2122 = n2120 & n2121;
  assign n2123 = ~n81 & n106;
  assign n2124 = ~n125 & ~n2123;
  assign n2125 = n2122 & n2124;
  assign n2126 = ~n233 & ~n460;
  assign n2127 = ~n824 & n2126;
  assign n2128 = n675 & n2127;
  assign n2129 = n2125 & n2128;
  assign n2130 = n2118 & n2129;
  assign n2131 = n202 & n2130;
  assign n2104 = n1820 ^ n1259;
  assign n2105 = n1842 ^ n1259;
  assign n2106 = n2105 ^ n1833;
  assign n2107 = ~n2104 & n2106;
  assign n2108 = n2107 ^ n1833;
  assign n2109 = n2108 ^ n1834;
  assign n2132 = n2131 ^ n2109;
  assign n2135 = n110 & ~n304;
  assign n2136 = ~n314 & ~n2135;
  assign n2137 = ~n514 & n2136;
  assign n2138 = n2076 & n2137;
  assign n2139 = n872 & n1924;
  assign n2140 = n1962 & n2139;
  assign n2141 = n2138 & n2140;
  assign n2142 = n641 & n2116;
  assign n2143 = ~n236 & ~n2031;
  assign n2144 = ~n267 & ~n2143;
  assign n2145 = n2142 & n2144;
  assign n2146 = ~n110 & n427;
  assign n2147 = ~n86 & n163;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = ~n215 & ~n2148;
  assign n2150 = n106 & ~n999;
  assign n2151 = n60 & ~n855;
  assign n2152 = ~n2150 & ~n2151;
  assign n2153 = ~n179 & n2152;
  assign n2154 = n2149 & n2153;
  assign n2155 = n219 & n1072;
  assign n2156 = ~n186 & ~n2155;
  assign n2157 = ~n93 & n2156;
  assign n2158 = n906 & n2157;
  assign n2159 = n2154 & n2158;
  assign n2160 = n2145 & n2159;
  assign n2161 = n2141 & n2160;
  assign n2162 = n735 & n2161;
  assign n2133 = n1831 ^ n1828;
  assign n2134 = n2133 ^ n2104;
  assign n2163 = n2162 ^ n2134;
  assign n2174 = n109 & ~n115;
  assign n2175 = n1963 & ~n2174;
  assign n2176 = n1923 & n2175;
  assign n2177 = ~n131 & ~n521;
  assign n2178 = n86 & ~n828;
  assign n2179 = ~n434 & ~n2178;
  assign n2180 = n2177 & n2179;
  assign n2181 = ~n59 & n159;
  assign n2182 = ~n45 & n136;
  assign n2183 = ~n55 & n2182;
  assign n2184 = ~n2181 & ~n2183;
  assign n2185 = n45 & n270;
  assign n2186 = n2184 & ~n2185;
  assign n2187 = n94 & ~n166;
  assign n2188 = ~n2186 & ~n2187;
  assign n2189 = n2180 & n2188;
  assign n2190 = n2176 & n2189;
  assign n253 = ~n251 & ~n252;
  assign n2191 = ~n676 & ~n721;
  assign n2192 = ~n168 & n2191;
  assign n2193 = n253 & n2192;
  assign n2194 = ~n436 & ~n472;
  assign n2195 = n2115 & n2194;
  assign n2196 = n2193 & n2195;
  assign n2197 = ~n242 & ~n2123;
  assign n2198 = n60 & ~n512;
  assign n2199 = n2197 & ~n2198;
  assign n2200 = n658 & n2199;
  assign n2201 = n2196 & n2200;
  assign n2202 = n2190 & n2201;
  assign n2203 = n2084 & n2202;
  assign n2172 = n1793 ^ n1790;
  assign n2164 = n1769 ^ n1766;
  assign n2173 = n2172 ^ n2164;
  assign n2204 = n2203 ^ n2173;
  assign n2205 = n1753 ^ n1750;
  assign n2209 = ~n1759 & n1760;
  assign n2206 = n1762 ^ n1757;
  assign n2207 = n2206 ^ n1757;
  assign n2208 = n2207 ^ n1753;
  assign n2210 = n2209 ^ n2208;
  assign n2211 = n2205 & n2210;
  assign n2212 = n2211 ^ n2209;
  assign n2213 = n2212 ^ n1745;
  assign n2214 = ~n61 & ~n1019;
  assign n2215 = n94 & ~n159;
  assign n2216 = n59 & ~n655;
  assign n2217 = ~n2215 & ~n2216;
  assign n2218 = ~n183 & n2217;
  assign n2219 = n703 & n2218;
  assign n2220 = n417 & n1029;
  assign n2221 = n2219 & n2220;
  assign n2222 = n734 & n869;
  assign n2223 = n2221 & n2222;
  assign n2224 = n2141 & n2223;
  assign n2225 = n1915 & n2224;
  assign n2226 = ~n2214 & n2225;
  assign n2227 = n2213 & n2226;
  assign n2228 = n2227 ^ n2203;
  assign n2229 = ~n2204 & ~n2228;
  assign n2230 = n2229 ^ n2173;
  assign n2166 = n1793 ^ n1789;
  assign n2167 = ~n1790 & n2166;
  assign n2165 = n1815 ^ n1769;
  assign n2168 = n2167 ^ n2165;
  assign n2169 = ~n2164 & ~n2168;
  assign n2170 = n2169 ^ n2167;
  assign n2171 = n2170 ^ n1808;
  assign n2231 = n2230 ^ n2171;
  assign n2232 = ~n183 & n361;
  assign n2233 = ~n274 & ~n326;
  assign n2234 = ~n472 & ~n712;
  assign n2235 = n2233 & n2234;
  assign n2236 = n2232 & n2235;
  assign n2238 = n896 & n2237;
  assign n2239 = n2236 & n2238;
  assign n2240 = n2154 & n2239;
  assign n245 = ~n241 & n244;
  assign n246 = n240 & n245;
  assign n2241 = n246 & n487;
  assign n2242 = n2240 & n2241;
  assign n2243 = n1999 & n2115;
  assign n2244 = ~n403 & ~n507;
  assign n2245 = ~n923 & n2244;
  assign n2246 = n161 & n2245;
  assign n2247 = n2243 & n2246;
  assign n2248 = ~n539 & ~n1043;
  assign n2250 = ~n271 & n2249;
  assign n2251 = n2248 & n2250;
  assign n2252 = n2247 & n2251;
  assign n2253 = n189 & n2091;
  assign n2254 = n2252 & n2253;
  assign n2255 = n2242 & n2254;
  assign n2256 = n2255 ^ n2230;
  assign n2257 = ~n2231 & n2256;
  assign n2258 = n2257 ^ n2171;
  assign n2259 = n2258 ^ n2134;
  assign n2260 = ~n2163 & n2259;
  assign n2261 = n2260 ^ n2258;
  assign n2262 = n2261 ^ n2131;
  assign n2263 = n2132 & ~n2262;
  assign n2264 = n2263 ^ n2109;
  assign n2265 = n2264 ^ n2102;
  assign n2266 = ~n2103 & n2265;
  assign n2267 = n2266 ^ n2264;
  assign n2268 = n2267 ^ n2074;
  assign n2269 = n2075 & ~n2268;
  assign n2270 = n2269 ^ n2267;
  assign n2271 = n2270 ^ n1990;
  assign n2272 = ~n2023 & n2271;
  assign n2273 = n2272 ^ n2270;
  assign n2274 = n2273 ^ n1947;
  assign n2275 = n1987 & ~n2274;
  assign n2276 = n2275 ^ n2273;
  assign n1941 = n1896 ^ n802;
  assign n2277 = n2276 ^ n1941;
  assign n2278 = ~n235 & ~n507;
  assign n2279 = ~n426 & n2278;
  assign n2280 = n230 & ~n444;
  assign n2281 = n2279 & n2280;
  assign n2282 = n219 & ~n1085;
  assign n2283 = ~n277 & ~n721;
  assign n2284 = ~n2282 & n2283;
  assign n2285 = n415 & n2284;
  assign n2286 = n2281 & n2285;
  assign n2287 = n480 & n648;
  assign n2288 = n732 & n2287;
  assign n2289 = n393 & n2288;
  assign n2290 = n2286 & n2289;
  assign n2291 = n1032 & n2290;
  assign n2292 = ~n521 & n943;
  assign n2293 = n2291 & n2292;
  assign n2294 = n2293 ^ n1941;
  assign n2295 = n2277 & ~n2294;
  assign n2296 = n2295 ^ n2276;
  assign n2297 = n2296 ^ n1900;
  assign n2298 = ~n1940 & n2297;
  assign n2299 = n2298 ^ n2296;
  assign n247 = n224 & n246;
  assign n254 = n250 & n253;
  assign n261 = ~n111 & ~n260;
  assign n262 = n259 & n261;
  assign n263 = n254 & n262;
  assign n265 = n110 & ~n236;
  assign n266 = ~n264 & ~n265;
  assign n272 = ~n267 & ~n271;
  assign n273 = n266 & n272;
  assign n276 = ~n274 & ~n275;
  assign n279 = ~n277 & ~n278;
  assign n280 = n276 & n279;
  assign n281 = n273 & n280;
  assign n282 = n263 & n281;
  assign n283 = n247 & n282;
  assign n284 = n202 & n283;
  assign n2300 = n2299 ^ n284;
  assign n2301 = n572 & n611;
  assign n2302 = ~n565 & ~n2301;
  assign n2303 = ~n318 & n2302;
  assign n2304 = ~n610 & ~n2303;
  assign n2310 = n609 & ~n2304;
  assign n2305 = ~n572 & ~n611;
  assign n2306 = ~n318 & n2305;
  assign n2311 = n546 & ~n565;
  assign n2312 = n2306 & n2311;
  assign n2313 = ~n2310 & ~n2312;
  assign n2314 = n1899 & ~n2313;
  assign n2404 = n2314 ^ n284;
  assign n2405 = n2300 & ~n2404;
  assign n2406 = n2405 ^ n2299;
  assign n3064 = n2403 & n2406;
  assign n3071 = ~n197 & n1913;
  assign n3072 = n1044 & n2177;
  assign n3073 = n3071 & n3072;
  assign n3074 = ~n314 & ~n491;
  assign n3075 = ~n298 & n3074;
  assign n3076 = n3073 & n3075;
  assign n3077 = n3070 & n3076;
  assign n3078 = n686 & n3077;
  assign n3079 = ~n248 & ~n271;
  assign n3080 = ~n414 & n3079;
  assign n3081 = ~n93 & ~n1049;
  assign n3082 = ~n687 & n2044;
  assign n3083 = n3081 & n3082;
  assign n3084 = n3080 & n3083;
  assign n3085 = n101 & n141;
  assign n3086 = ~n1005 & ~n3085;
  assign n3087 = n3084 & ~n3086;
  assign n3088 = ~n461 & ~n887;
  assign n3089 = n60 & ~n999;
  assign n3090 = ~n319 & ~n3089;
  assign n3091 = n3088 & n3090;
  assign n3092 = n1935 & n3091;
  assign n3093 = n3087 & n3092;
  assign n3094 = n725 & n3093;
  assign n3095 = n3078 & n3094;
  assign n3096 = n3064 & n3095;
  assign n3115 = n3063 & n3096;
  assign n3630 = n3114 & n3115;
  assign n3631 = ~n105 & n3102;
  assign n3632 = n71 & n236;
  assign n3633 = n109 & ~n3632;
  assign n3634 = ~n314 & ~n3633;
  assign n3635 = ~n682 & n3634;
  assign n3636 = n256 & n306;
  assign n3637 = ~n84 & n3636;
  assign n3638 = n55 & ~n3637;
  assign n3639 = n2124 & ~n3638;
  assign n3640 = n3635 & n3639;
  assign n3641 = n313 & n3640;
  assign n3642 = n3631 & n3641;
  assign n3643 = ~n3630 & ~n3642;
  assign n3644 = n3267 & n3643;
  assign n3116 = n3115 ^ n3114;
  assign n3188 = ~x0 & x1;
  assign n3645 = ~n3116 & n3188;
  assign n3097 = n3096 ^ n3063;
  assign n3249 = ~x0 & n2322;
  assign n3646 = ~n3097 & n3249;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n3644 & n3647;
  assign n3649 = n2323 & ~n3648;
  assign n3179 = x1 & ~x2;
  assign n3180 = x0 & x22;
  assign n3181 = n3179 & n3180;
  assign n2324 = ~n26 & ~n2323;
  assign n3205 = x22 ^ x1;
  assign n3206 = x0 & n3205;
  assign n3657 = n2324 & ~n3206;
  assign n3658 = n3648 & n3657;
  assign n3659 = ~n3181 & ~n3658;
  assign n2307 = n2304 & ~n2306;
  assign n2308 = n2307 ^ n1899;
  assign n2309 = n615 & n2308;
  assign n2315 = n2314 ^ n2309;
  assign n2316 = ~n2300 & ~n2315;
  assign n2317 = n2316 ^ n2314;
  assign n2320 = n2296 ^ n1940;
  assign n2342 = n2273 ^ n1987;
  assign n2343 = n2270 ^ n2023;
  assign n2344 = n2267 ^ n2075;
  assign n2345 = n2264 ^ n2103;
  assign n2346 = n2261 ^ n2132;
  assign n2347 = n2258 ^ n2163;
  assign n2348 = n2255 ^ n2171;
  assign n2349 = n2348 ^ n2230;
  assign n2350 = n2227 ^ n2204;
  assign n2351 = n2349 & n2350;
  assign n2352 = n2347 & ~n2351;
  assign n2353 = ~n2346 & ~n2352;
  assign n2354 = n2345 & ~n2353;
  assign n2355 = n2344 & ~n2354;
  assign n2356 = n2343 & ~n2355;
  assign n2357 = n2342 & ~n2356;
  assign n2358 = n2293 ^ n1940;
  assign n2359 = n2293 ^ n2276;
  assign n2360 = n2293 ^ n2277;
  assign n2361 = ~n2293 & n2360;
  assign n2362 = n2361 ^ n2293;
  assign n2363 = ~n2359 & ~n2362;
  assign n2364 = n2363 ^ n2361;
  assign n2365 = n2364 ^ n2293;
  assign n2366 = n2365 ^ n2277;
  assign n2367 = ~n2358 & n2366;
  assign n2368 = n2367 ^ n1940;
  assign n2369 = ~n2357 & ~n2368;
  assign n2370 = ~n2320 & ~n2369;
  assign n3119 = ~n2317 & ~n2370;
  assign n3120 = ~n2403 & ~n2406;
  assign n3121 = ~n3119 & n3120;
  assign n3122 = n3095 & ~n3121;
  assign n3123 = n3064 & n3119;
  assign n3124 = ~n3063 & ~n3123;
  assign n3125 = ~n3122 & n3124;
  assign n3650 = n3114 & ~n3115;
  assign n3651 = ~n3125 & n3650;
  assign n3126 = ~n3064 & ~n3095;
  assign n2371 = n2226 ^ n2213;
  assign n2372 = n2350 & ~n2371;
  assign n2373 = ~n2349 & ~n2372;
  assign n2374 = ~n2347 & ~n2373;
  assign n2375 = n2346 & ~n2374;
  assign n2376 = ~n2345 & ~n2375;
  assign n2377 = ~n2344 & ~n2376;
  assign n2378 = ~n2343 & ~n2377;
  assign n2379 = ~n2342 & ~n2378;
  assign n2380 = ~n2360 & ~n2379;
  assign n2381 = n2320 & ~n2380;
  assign n3131 = ~n284 & ~n2299;
  assign n3132 = ~n2309 & n3131;
  assign n3133 = ~n2381 & n3132;
  assign n3127 = n284 & n2299;
  assign n3128 = n2309 & n3127;
  assign n3129 = n2381 & n2406;
  assign n3130 = ~n3128 & ~n3129;
  assign n3134 = n3133 ^ n3130;
  assign n3135 = n3134 ^ n3130;
  assign n3136 = n3130 ^ n2406;
  assign n3137 = n3136 ^ n3130;
  assign n3138 = ~n3135 & ~n3137;
  assign n3139 = n3138 ^ n3130;
  assign n3140 = n2403 & ~n3139;
  assign n3141 = n3140 ^ n3130;
  assign n3142 = n3126 & n3141;
  assign n3143 = n3063 & ~n3142;
  assign n3652 = n3143 ^ n3115;
  assign n3653 = n3114 & ~n3652;
  assign n3654 = n3653 ^ n3143;
  assign n3655 = ~n3651 & n3654;
  assign n3656 = n3655 ^ n3643;
  assign n3660 = n3659 ^ n3656;
  assign n3661 = n3660 ^ n3659;
  assign n2325 = x0 & ~x22;
  assign n2326 = x2 & n2325;
  assign n2327 = n2324 & ~n2326;
  assign n3662 = n2327 & n3648;
  assign n3663 = n3662 ^ n3659;
  assign n3664 = ~n3661 & ~n3663;
  assign n3665 = n3664 ^ n3659;
  assign n3666 = ~n3649 & n3665;
  assign n2590 = n596 & ~n2371;
  assign n2451 = n618 ^ n595;
  assign n2483 = n2204 & n2371;
  assign n2591 = n2451 & n2483;
  assign n2592 = n2591 ^ n2349;
  assign n2593 = n1108 & n2592;
  assign n2449 = n621 & ~n1108;
  assign n2594 = n2350 & n2449;
  assign n2453 = ~n620 & ~n812;
  assign n2452 = n620 & n812;
  assign n2454 = n2453 ^ n2452;
  assign n2455 = n2452 ^ n618;
  assign n2456 = n2455 ^ n2452;
  assign n2457 = n2454 & ~n2456;
  assign n2458 = n2457 ^ n2452;
  assign n2459 = n2451 & n2458;
  assign n2595 = ~n2371 & n2459;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = ~n2593 & n2596;
  assign n2598 = n618 & ~n2371;
  assign n2599 = n2453 & ~n2598;
  assign n2600 = n2452 ^ n2371;
  assign n2601 = n2452 ^ n2204;
  assign n2602 = n2601 ^ n2204;
  assign n2603 = n2204 ^ n618;
  assign n2604 = n2602 & n2603;
  assign n2605 = n2604 ^ n2204;
  assign n2606 = n2600 & n2605;
  assign n2607 = n2606 ^ n2371;
  assign n2608 = ~n2599 & ~n2607;
  assign n2609 = n595 & ~n2608;
  assign n2610 = n2597 & n2609;
  assign n2611 = ~n2590 & ~n2610;
  assign n2612 = n2349 & n2449;
  assign n2613 = n2350 & n2459;
  assign n2614 = ~n2612 & ~n2613;
  assign n2500 = ~n2351 & ~n2373;
  assign n2615 = n618 & n2500;
  assign n2616 = n2615 ^ n2347;
  assign n2617 = n1108 & ~n2616;
  assign n2618 = n2617 ^ n595;
  assign n2619 = n2618 ^ n2617;
  assign n2620 = ~n618 & n2500;
  assign n2621 = n2620 ^ n2347;
  assign n2622 = n1108 & ~n2621;
  assign n2623 = n2622 ^ n2617;
  assign n2624 = n2619 & n2623;
  assign n2625 = n2624 ^ n2617;
  assign n2626 = n2614 & ~n2625;
  assign n2627 = n2626 ^ n595;
  assign n2628 = ~n2611 & ~n2627;
  assign n2580 = n2371 ^ n2350;
  assign n2581 = n2580 ^ n2350;
  assign n2582 = n2350 ^ n579;
  assign n2583 = n2582 ^ n2350;
  assign n2584 = ~n2581 & n2583;
  assign n2585 = n2584 ^ n2350;
  assign n2586 = ~n596 & n2585;
  assign n2587 = n2586 ^ n2350;
  assign n2474 = ~n572 & ~n2371;
  assign n2588 = n2587 ^ n2474;
  assign n2560 = ~n2352 & ~n2374;
  assign n2561 = n1108 & ~n2346;
  assign n2562 = ~n2560 & n2561;
  assign n2563 = ~n2347 & n2449;
  assign n2564 = n2349 & n2459;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = ~n2562 & n2565;
  assign n2567 = ~n595 & ~n2566;
  assign n2568 = n1108 & n2560;
  assign n2569 = n2346 ^ n618;
  assign n2570 = n2569 ^ n2561;
  assign n2571 = n2570 ^ n2569;
  assign n2572 = n595 & n2565;
  assign n2573 = n2572 ^ n2569;
  assign n2574 = n2573 ^ n2569;
  assign n2575 = ~n2571 & n2574;
  assign n2576 = n2575 ^ n2569;
  assign n2577 = ~n2568 & ~n2576;
  assign n2578 = n2577 ^ n2569;
  assign n2579 = ~n2567 & n2578;
  assign n2589 = n2588 ^ n2579;
  assign n2673 = n2628 ^ n2589;
  assign n2656 = ~n2355 & ~n2377;
  assign n2657 = ~n2343 & ~n2656;
  assign n2658 = n1451 & n2657;
  assign n2425 = ~n30 & ~n1100;
  assign n2424 = n30 & n1100;
  assign n2426 = n2425 ^ n2424;
  assign n2427 = n816 & n2426;
  assign n2428 = n2427 ^ n2425;
  assign n2659 = n2344 & n2428;
  assign n2430 = n2427 ^ n2424;
  assign n2431 = ~n817 & n2430;
  assign n2660 = ~n2345 & n2431;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2658 & n2661;
  assign n2663 = ~n812 & ~n2662;
  assign n2664 = n2343 & ~n2656;
  assign n2665 = n1451 & ~n2664;
  assign n2666 = n812 & n2661;
  assign n2667 = ~n2665 & n2666;
  assign n2668 = n1451 & n2656;
  assign n2669 = n2343 ^ n816;
  assign n2670 = n2668 & n2669;
  assign n2671 = ~n2667 & ~n2670;
  assign n2672 = ~n2663 & n2671;
  assign n2674 = n2673 ^ n2672;
  assign n2690 = n595 & n2614;
  assign n2691 = ~n2622 & n2690;
  assign n2692 = ~n2590 & n2691;
  assign n2689 = n2627 ^ n2590;
  assign n2693 = n2692 ^ n2689;
  assign n2694 = n2610 & n2693;
  assign n2695 = n2694 ^ n2689;
  assign n2445 = ~n2354 & ~n2376;
  assign n2463 = n2344 & ~n2445;
  assign n2675 = n1451 & n2463;
  assign n2676 = ~n2345 & n2428;
  assign n2677 = ~n2346 & n2431;
  assign n2678 = ~n2676 & ~n2677;
  assign n2679 = ~n2675 & n2678;
  assign n2680 = ~n812 & ~n2679;
  assign n2466 = ~n2344 & ~n2445;
  assign n2681 = n1451 & ~n2466;
  assign n2682 = n812 & n2678;
  assign n2683 = ~n2681 & n2682;
  assign n2684 = n1451 & n2445;
  assign n2685 = n2344 ^ n816;
  assign n2686 = n2684 & ~n2685;
  assign n2687 = ~n2683 & ~n2686;
  assign n2688 = ~n2680 & n2687;
  assign n2696 = n2695 ^ n2688;
  assign n2735 = n2350 ^ n620;
  assign n2736 = n2735 ^ n2350;
  assign n2737 = ~n2581 & n2736;
  assign n2738 = n2737 ^ n2350;
  assign n2739 = ~n1108 & n2738;
  assign n2740 = n2739 ^ n2350;
  assign n2741 = n2740 ^ n2598;
  assign n2699 = ~n817 & n2483;
  assign n2700 = n2699 ^ n2349;
  assign n2701 = n1451 & n2700;
  assign n2702 = n2350 & n2428;
  assign n2703 = ~n2371 & n2431;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~n2701 & n2704;
  assign n2706 = n1451 & n2350;
  assign n2707 = n2371 & ~n2706;
  assign n2708 = ~n2430 & ~n2707;
  assign n2709 = n812 & ~n2708;
  assign n2710 = n2705 & n2709;
  assign n2711 = n1108 & ~n2371;
  assign n2712 = ~n2710 & ~n2711;
  assign n2713 = n2349 & n2428;
  assign n2714 = n2350 & n2431;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = n2715 ^ n812;
  assign n2717 = n2347 & ~n2500;
  assign n2718 = n1451 & ~n2717;
  assign n2719 = n2718 ^ n2715;
  assign n2720 = ~n812 & ~n2500;
  assign n2721 = n1451 & ~n2720;
  assign n2722 = n816 & n2500;
  assign n2723 = n2722 ^ n2347;
  assign n2724 = n2721 & ~n2723;
  assign n2725 = n2724 ^ n2715;
  assign n2726 = n2715 & ~n2725;
  assign n2727 = n2726 ^ n2715;
  assign n2728 = n2719 & n2727;
  assign n2729 = n2728 ^ n2726;
  assign n2730 = n2729 ^ n2715;
  assign n2731 = n2730 ^ n2724;
  assign n2732 = n2716 & ~n2731;
  assign n2733 = n2732 ^ n2724;
  assign n2734 = ~n2712 & ~n2733;
  assign n2742 = n2741 ^ n2734;
  assign n2743 = n2560 ^ n2346;
  assign n2744 = ~n816 & n1451;
  assign n2745 = ~n2743 & n2744;
  assign n2746 = n812 & ~n816;
  assign n2747 = ~n2347 & n2428;
  assign n2748 = n2349 & n2431;
  assign n2749 = ~n2747 & ~n2748;
  assign n2750 = ~n2746 & n2749;
  assign n2751 = n816 & n1451;
  assign n2752 = ~n2346 & n2751;
  assign n2753 = n2750 & ~n2752;
  assign n2754 = ~n2745 & n2753;
  assign n2755 = n2346 & n2749;
  assign n2756 = n812 & ~n2755;
  assign n2757 = ~n2754 & ~n2756;
  assign n2758 = n1451 & ~n2743;
  assign n2759 = n812 & ~n2744;
  assign n2760 = n2749 & n2759;
  assign n2761 = ~n2758 & n2760;
  assign n2762 = ~n2757 & ~n2761;
  assign n2763 = n2762 ^ n2741;
  assign n2764 = n2742 & n2763;
  assign n2765 = n2764 ^ n2734;
  assign n2697 = n595 & n2608;
  assign n2698 = n2697 ^ n2597;
  assign n2766 = n2765 ^ n2698;
  assign n2525 = ~n2353 & ~n2375;
  assign n2767 = ~n2345 & ~n2525;
  assign n2768 = n1451 & n2767;
  assign n2769 = ~n2346 & n2428;
  assign n2770 = ~n2347 & n2431;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = ~n2768 & n2771;
  assign n2773 = n812 & ~n2772;
  assign n2541 = n2345 & ~n2525;
  assign n2774 = n1451 & ~n2541;
  assign n2775 = ~n812 & n2771;
  assign n2776 = ~n2774 & n2775;
  assign n2777 = n1451 & n2525;
  assign n2778 = n2345 ^ n816;
  assign n2779 = n2777 & ~n2778;
  assign n2780 = ~n2776 & ~n2779;
  assign n2781 = ~n2773 & n2780;
  assign n2782 = n2781 ^ n2698;
  assign n2783 = n2766 & ~n2782;
  assign n2784 = n2783 ^ n2781;
  assign n2785 = n2784 ^ n2688;
  assign n2786 = ~n2696 & ~n2785;
  assign n2787 = n2786 ^ n2784;
  assign n2788 = n2787 ^ n2672;
  assign n2789 = ~n2674 & ~n2788;
  assign n2790 = n2789 ^ n2787;
  assign n2629 = n2628 ^ n2588;
  assign n2630 = ~n2589 & ~n2629;
  assign n2631 = n2630 ^ n2579;
  assign n2473 = ~n2204 & n2371;
  assign n2475 = ~n565 & n611;
  assign n2476 = ~n2474 & n2475;
  assign n2477 = ~n2473 & ~n2476;
  assign n2478 = n579 & n595;
  assign n2479 = n572 & n2478;
  assign n2480 = ~n2371 & n2479;
  assign n2481 = n2480 ^ n2478;
  assign n2482 = n2477 & ~n2481;
  assign n2557 = ~n565 & n2482;
  assign n2484 = n573 & n2483;
  assign n2485 = n2484 ^ n2349;
  assign n2486 = n596 & n2485;
  assign n2487 = ~n572 & n611;
  assign n2488 = ~n2479 & ~n2487;
  assign n2489 = n2350 & ~n2488;
  assign n2490 = n565 & n2478;
  assign n2491 = ~n2475 & ~n2490;
  assign n2492 = n573 & ~n2491;
  assign n2493 = ~n2371 & n2492;
  assign n2494 = ~n2489 & ~n2493;
  assign n2495 = ~n2486 & n2494;
  assign n2558 = n2557 ^ n2495;
  assign n2526 = ~n618 & n2525;
  assign n2527 = ~n2345 & ~n2526;
  assign n2528 = ~n2346 & n2449;
  assign n2529 = ~n2347 & n2459;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = n2530 ^ n1108;
  assign n2532 = n2531 ^ n1108;
  assign n2533 = n2525 ^ n1108;
  assign n2534 = n2533 ^ n1108;
  assign n2535 = n2532 & n2534;
  assign n2536 = n2535 ^ n1108;
  assign n2537 = ~n595 & n2536;
  assign n2538 = n2537 ^ n1108;
  assign n2539 = n2527 & n2538;
  assign n2540 = n2530 ^ n595;
  assign n2542 = n1108 & ~n2541;
  assign n2543 = n2542 ^ n595;
  assign n2544 = ~n618 & n1108;
  assign n2545 = n2345 & n2544;
  assign n2546 = n2525 & n2545;
  assign n2547 = n2546 ^ n595;
  assign n2548 = ~n595 & n2547;
  assign n2549 = n2548 ^ n595;
  assign n2550 = ~n2543 & ~n2549;
  assign n2551 = n2550 ^ n2548;
  assign n2552 = n2551 ^ n595;
  assign n2553 = n2552 ^ n2546;
  assign n2554 = n2540 & n2553;
  assign n2555 = n2554 ^ n2546;
  assign n2556 = ~n2539 & ~n2555;
  assign n2559 = n2558 ^ n2556;
  assign n2654 = n2631 ^ n2559;
  assign n2637 = ~n2356 & ~n2378;
  assign n2638 = n2342 & ~n2637;
  assign n2639 = n1451 & n2638;
  assign n2640 = ~n2343 & n2428;
  assign n2641 = n2344 & n2431;
  assign n2642 = ~n2640 & ~n2641;
  assign n2643 = ~n2639 & n2642;
  assign n2644 = n812 & ~n2643;
  assign n2645 = ~n2342 & ~n2637;
  assign n2646 = n1451 & ~n2645;
  assign n2647 = ~n812 & n2642;
  assign n2648 = ~n2646 & n2647;
  assign n2649 = n1451 & n2637;
  assign n2650 = n2342 ^ n816;
  assign n2651 = n2649 & n2650;
  assign n2652 = ~n2648 & ~n2651;
  assign n2653 = ~n2644 & n2652;
  assign n2655 = n2654 ^ n2653;
  assign n2822 = n2790 ^ n2655;
  assign n2385 = n2327 ^ n1323;
  assign n2382 = ~n2370 & ~n2381;
  assign n2795 = n32 ^ n30;
  assign n2796 = n2382 & n2795;
  assign n2797 = n2796 ^ n30;
  assign n2798 = n2797 ^ n2317;
  assign n2799 = n2385 & ~n2798;
  assign n2333 = n1323 & n2327;
  assign n2334 = ~n32 & n2333;
  assign n2328 = ~n1323 & ~n2327;
  assign n2802 = n32 & n2328;
  assign n2803 = ~n2334 & ~n2802;
  assign n2804 = n30 & ~n2803;
  assign n2800 = ~n2328 & ~n2334;
  assign n2801 = ~n30 & ~n2800;
  assign n2805 = n2804 ^ n2801;
  assign n2806 = ~n2320 & n2805;
  assign n2807 = n2806 ^ n2801;
  assign n2336 = ~n30 & n32;
  assign n2337 = n2333 & n2336;
  assign n2329 = ~n32 & n2328;
  assign n2808 = n2337 ^ n2329;
  assign n2809 = n2808 ^ n2329;
  assign n2810 = n2809 ^ n2329;
  assign n2811 = n2360 ^ n2329;
  assign n2812 = n2811 ^ n2329;
  assign n2813 = n2810 & n2812;
  assign n2814 = n2813 ^ n2329;
  assign n2815 = ~n30 & n2329;
  assign n2816 = n2815 ^ n2807;
  assign n2817 = n2814 & ~n2816;
  assign n2818 = n2817 ^ n2815;
  assign n2819 = ~n2807 & n2818;
  assign n2820 = n2819 ^ n2807;
  assign n2821 = ~n2799 & ~n2820;
  assign n2823 = n2822 ^ n2821;
  assign n2825 = n2360 ^ n2342;
  assign n2826 = n2825 ^ n2360;
  assign n2827 = n2360 ^ n30;
  assign n2828 = n2827 ^ n2360;
  assign n2829 = n2826 & n2828;
  assign n2830 = n2829 ^ n2360;
  assign n2831 = ~n32 & ~n2830;
  assign n2832 = n2831 ^ n2360;
  assign n2833 = n2328 & ~n2832;
  assign n2834 = n2334 & ~n2360;
  assign n2835 = n2337 & n2342;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = ~n2833 & n2836;
  assign n2838 = n2837 ^ n30;
  assign n2839 = n2379 ^ n2357;
  assign n2840 = n2360 & n2839;
  assign n2841 = n2840 ^ n2379;
  assign n2842 = n2320 & ~n2841;
  assign n2843 = n2385 & ~n2842;
  assign n2844 = n2843 ^ n30;
  assign n2845 = ~n30 & n2385;
  assign n2846 = ~n2320 & ~n2841;
  assign n2847 = n2845 & n2846;
  assign n2848 = n2320 ^ n32;
  assign n2849 = n2385 & n2841;
  assign n2850 = ~n2848 & n2849;
  assign n2851 = ~n2847 & ~n2850;
  assign n2852 = n2851 ^ n30;
  assign n2853 = n30 & n2852;
  assign n2854 = n2853 ^ n30;
  assign n2855 = n2844 & n2854;
  assign n2856 = n2855 ^ n2853;
  assign n2857 = n2856 ^ n30;
  assign n2858 = n2857 ^ n2851;
  assign n2859 = ~n2838 & n2858;
  assign n2860 = n2859 ^ n2851;
  assign n2824 = n2787 ^ n2674;
  assign n2861 = n2860 ^ n2824;
  assign n2880 = n2784 ^ n2696;
  assign n2412 = n30 & n2385;
  assign n2421 = ~n2357 & ~n2379;
  assign n2422 = ~n2360 & ~n2421;
  assign n2862 = n2412 & n2422;
  assign n2863 = n2342 & ~n2803;
  assign n2864 = n1323 ^ n32;
  assign n2865 = n2327 ^ n32;
  assign n2866 = ~n2864 & ~n2865;
  assign n2867 = n2795 & n2866;
  assign n2868 = ~n2343 & n2867;
  assign n2869 = ~n2863 & ~n2868;
  assign n2870 = n30 & ~n2869;
  assign n2871 = ~n2862 & ~n2870;
  assign n2872 = n2360 ^ n32;
  assign n2873 = n2385 & n2421;
  assign n2874 = n2872 & n2873;
  assign n2875 = n2871 & ~n2874;
  assign n2436 = n2360 & ~n2421;
  assign n2876 = n2385 & ~n2436;
  assign n2877 = ~n30 & n2869;
  assign n2878 = ~n2876 & n2877;
  assign n2879 = n2875 & ~n2878;
  assign n2881 = n2880 ^ n2879;
  assign n2896 = n2781 ^ n2766;
  assign n2882 = n2385 & ~n2645;
  assign n2883 = ~n2343 & ~n2803;
  assign n2884 = n2344 & n2867;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = n30 & n2885;
  assign n2887 = ~n2882 & n2886;
  assign n2888 = n2385 & n2637;
  assign n2889 = n2342 ^ n32;
  assign n2890 = n2888 & n2889;
  assign n2891 = ~n2887 & ~n2890;
  assign n2892 = n2638 & n2845;
  assign n2893 = ~n30 & ~n2885;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = n2891 & n2894;
  assign n2897 = n2896 ^ n2895;
  assign n2918 = n2762 ^ n2742;
  assign n2898 = n2385 & n2656;
  assign n2899 = n2343 ^ n32;
  assign n2900 = n2898 & n2899;
  assign n2901 = n2344 & ~n2803;
  assign n2902 = ~n2345 & n2867;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n2903 ^ n30;
  assign n2905 = n2385 & ~n2664;
  assign n2906 = n2905 ^ n2903;
  assign n2907 = n2412 & n2657;
  assign n2908 = n2907 ^ n2905;
  assign n2909 = n2905 & ~n2908;
  assign n2910 = n2909 ^ n2905;
  assign n2911 = n2906 & n2910;
  assign n2912 = n2911 ^ n2909;
  assign n2913 = n2912 ^ n2905;
  assign n2914 = n2913 ^ n2907;
  assign n2915 = n2904 & ~n2914;
  assign n2916 = n2915 ^ n2907;
  assign n2917 = ~n2900 & ~n2916;
  assign n2919 = n2918 ^ n2917;
  assign n2950 = n2733 ^ n2712;
  assign n2951 = n2710 & n2711;
  assign n2952 = ~n2950 & ~n2951;
  assign n2920 = n32 & n2445;
  assign n2921 = n2344 & ~n2920;
  assign n2922 = ~n2345 & ~n2803;
  assign n2923 = ~n2346 & n2867;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n2924 ^ n2385;
  assign n2926 = n2925 ^ n2385;
  assign n2927 = n2445 ^ n2385;
  assign n2928 = n2927 ^ n2385;
  assign n2929 = n2926 & n2928;
  assign n2930 = n2929 ^ n2385;
  assign n2931 = n30 & n2930;
  assign n2932 = n2931 ^ n2385;
  assign n2933 = n2921 & n2932;
  assign n2934 = n2924 ^ n30;
  assign n2935 = n2385 & ~n2466;
  assign n2936 = n2935 ^ n30;
  assign n2937 = ~n2344 & n2445;
  assign n2938 = n32 & n2385;
  assign n2939 = n2937 & n2938;
  assign n2940 = n2939 ^ n30;
  assign n2941 = n30 & ~n2940;
  assign n2942 = n2941 ^ n30;
  assign n2943 = n2936 & n2942;
  assign n2944 = n2943 ^ n2941;
  assign n2945 = n2944 ^ n30;
  assign n2946 = n2945 ^ n2939;
  assign n2947 = ~n2934 & ~n2946;
  assign n2948 = n2947 ^ n2939;
  assign n2949 = ~n2933 & ~n2948;
  assign n2953 = n2952 ^ n2949;
  assign n2968 = n812 & n2708;
  assign n2969 = n2968 ^ n2705;
  assign n2954 = n2767 & n2845;
  assign n2955 = ~n2346 & ~n2803;
  assign n2956 = ~n2347 & n2867;
  assign n2957 = ~n2955 & ~n2956;
  assign n2958 = ~n30 & ~n2957;
  assign n2959 = ~n2954 & ~n2958;
  assign n2960 = n2345 ^ n32;
  assign n2961 = n2385 & n2525;
  assign n2962 = ~n2960 & n2961;
  assign n2963 = n2959 & ~n2962;
  assign n2964 = n2385 & ~n2541;
  assign n2965 = n30 & n2957;
  assign n2966 = ~n2964 & n2965;
  assign n2967 = n2963 & ~n2966;
  assign n2970 = n2969 ^ n2967;
  assign n3006 = n2424 ^ n816;
  assign n3007 = ~n2371 & ~n3006;
  assign n3008 = n3007 ^ n2706;
  assign n2971 = n2500 & n2795;
  assign n2972 = n2971 ^ n2347;
  assign n2973 = n2385 & ~n2972;
  assign n2974 = n2349 & ~n2803;
  assign n2975 = n2350 & n2867;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = ~n2973 & n2976;
  assign n2996 = ~n30 & n1100;
  assign n2997 = ~n2371 & n2996;
  assign n2978 = ~n2473 & ~n2866;
  assign n2979 = n30 & ~n2978;
  assign n33 = n30 & ~n32;
  assign n2982 = n2336 ^ n33;
  assign n2983 = n1323 & n2982;
  assign n2984 = n2983 ^ n33;
  assign n2985 = ~n2371 & n2984;
  assign n2980 = n2483 & n2795;
  assign n2981 = n2980 ^ n2349;
  assign n2986 = n2985 ^ n2981;
  assign n2987 = n2986 ^ n2981;
  assign n2988 = n2350 & n2864;
  assign n2989 = n2988 ^ n2981;
  assign n2990 = n2989 ^ n2981;
  assign n2991 = ~n2987 & ~n2990;
  assign n2992 = n2991 ^ n2981;
  assign n2993 = ~n2385 & ~n2992;
  assign n2994 = n2993 ^ n2981;
  assign n2995 = n2979 & ~n2994;
  assign n2998 = n2997 ^ n2995;
  assign n2999 = n2998 ^ n2997;
  assign n3000 = n1451 & ~n2371;
  assign n3001 = n3000 ^ n2997;
  assign n3002 = ~n2999 & ~n3001;
  assign n3003 = n3002 ^ n2997;
  assign n3004 = n2977 & ~n3003;
  assign n3005 = n3004 ^ n2997;
  assign n3009 = n3008 ^ n3005;
  assign n3013 = ~n2347 & n2864;
  assign n3014 = n2349 & n2984;
  assign n3015 = ~n3013 & ~n3014;
  assign n3016 = n3015 ^ n30;
  assign n3010 = n2560 & n2795;
  assign n3011 = n3010 ^ n30;
  assign n3012 = n3011 ^ n2346;
  assign n3017 = n3016 ^ n3012;
  assign n3018 = ~n2385 & n3017;
  assign n3019 = n3018 ^ n3012;
  assign n3020 = n3019 ^ n3008;
  assign n3021 = n3009 & n3020;
  assign n3022 = n3021 ^ n3005;
  assign n3023 = n3022 ^ n2969;
  assign n3024 = n2970 & n3023;
  assign n3025 = n3024 ^ n2967;
  assign n3026 = n3025 ^ n2952;
  assign n3027 = n2953 & ~n3026;
  assign n3028 = n3027 ^ n2949;
  assign n3029 = n3028 ^ n2918;
  assign n3030 = ~n2919 & ~n3029;
  assign n3031 = n3030 ^ n2917;
  assign n3032 = n3031 ^ n2896;
  assign n3033 = n2897 & n3032;
  assign n3034 = n3033 ^ n2895;
  assign n3035 = n3034 ^ n2880;
  assign n3036 = n2881 & n3035;
  assign n3037 = n3036 ^ n2879;
  assign n3038 = n3037 ^ n2860;
  assign n3039 = n2861 & ~n3038;
  assign n3040 = n3039 ^ n3037;
  assign n3041 = n3040 ^ n2822;
  assign n3042 = n2823 & ~n3041;
  assign n3043 = n3042 ^ n2821;
  assign n2791 = n2790 ^ n2654;
  assign n2792 = n2655 & ~n2791;
  assign n2793 = n2792 ^ n2653;
  assign n2632 = n2631 ^ n2558;
  assign n2633 = ~n2559 & ~n2632;
  assign n2634 = n2633 ^ n2556;
  assign n2496 = ~n2482 & n2495;
  assign n2497 = n2496 ^ n2371;
  assign n2498 = n2496 ^ n565;
  assign n2499 = n2498 ^ n565;
  assign n2501 = n573 & n2500;
  assign n2502 = n2501 ^ n2347;
  assign n2503 = n596 & n2502;
  assign n2507 = n565 & ~n572;
  assign n2508 = n2350 & n2507;
  assign n2509 = n2478 & ~n2508;
  assign n2504 = ~n565 & n572;
  assign n2505 = n2350 & n2504;
  assign n2506 = n611 & ~n2505;
  assign n2510 = n2509 ^ n2506;
  assign n2511 = n2349 ^ n572;
  assign n2512 = n2511 ^ n572;
  assign n2513 = n2509 ^ n572;
  assign n2514 = ~n2512 & ~n2513;
  assign n2515 = n2514 ^ n572;
  assign n2516 = n2510 & ~n2515;
  assign n2517 = n2516 ^ n2506;
  assign n2518 = ~n2503 & ~n2517;
  assign n2519 = n2518 ^ n565;
  assign n2520 = n2499 & n2519;
  assign n2521 = n2520 ^ n565;
  assign n2522 = n2497 & ~n2521;
  assign n2523 = n2522 ^ n2518;
  assign n2446 = n1108 & n2445;
  assign n2447 = n2344 ^ n618;
  assign n2448 = n2446 & ~n2447;
  assign n2450 = ~n2345 & n2449;
  assign n2460 = ~n2346 & n2459;
  assign n2461 = ~n2450 & ~n2460;
  assign n2462 = n2461 ^ n595;
  assign n2467 = n1108 & ~n2466;
  assign n2468 = ~n595 & n2467;
  assign n2464 = n595 & n1108;
  assign n2465 = n2463 & n2464;
  assign n2469 = n2468 ^ n2465;
  assign n2470 = n2462 & ~n2469;
  assign n2471 = n2470 ^ n2465;
  assign n2472 = ~n2448 & ~n2471;
  assign n2524 = n2523 ^ n2472;
  assign n2635 = n2634 ^ n2524;
  assign n2423 = n1451 & n2422;
  assign n2429 = n2342 & n2428;
  assign n2432 = ~n2343 & n2431;
  assign n2433 = ~n2429 & ~n2432;
  assign n2434 = ~n2423 & n2433;
  assign n2435 = n812 & ~n2434;
  assign n2437 = n1451 & ~n2436;
  assign n2438 = ~n812 & n2433;
  assign n2439 = ~n2437 & n2438;
  assign n2440 = n2360 ^ n816;
  assign n2441 = n1451 & n2421;
  assign n2442 = ~n2440 & n2441;
  assign n2443 = ~n2439 & ~n2442;
  assign n2444 = ~n2435 & n2443;
  assign n2636 = n2635 ^ n2444;
  assign n2794 = n2793 ^ n2636;
  assign n3044 = n3043 ^ n2794;
  assign n2318 = n32 & n2317;
  assign n2319 = ~n33 & ~n2318;
  assign n2330 = n2320 & n2329;
  assign n2331 = n2330 ^ n2328;
  assign n2332 = ~n2319 & n2331;
  assign n2335 = n2317 & n2334;
  assign n2338 = ~n2320 & n2337;
  assign n2339 = ~n2335 & ~n2338;
  assign n2340 = ~n2332 & n2339;
  assign n2341 = n30 & ~n2340;
  assign n2383 = n2320 ^ n2317;
  assign n2384 = ~n2382 & ~n2383;
  assign n2407 = n2406 ^ n2403;
  assign n2408 = n2407 ^ n32;
  assign n2409 = n2385 & n2408;
  assign n2410 = n2384 & n2409;
  assign n2411 = ~n2341 & ~n2410;
  assign n2413 = ~n2384 & ~n2407;
  assign n2414 = n2412 & n2413;
  assign n2415 = n2411 & ~n2414;
  assign n2416 = ~n30 & n2340;
  assign n2417 = ~n2384 & n2407;
  assign n2418 = n2385 & ~n2417;
  assign n2419 = n2416 & ~n2418;
  assign n2420 = n2415 & ~n2419;
  assign n3626 = n3043 ^ n2420;
  assign n3627 = ~n3044 & n3626;
  assign n3628 = n3627 ^ n2420;
  assign n3621 = n2793 ^ n2635;
  assign n3622 = n2636 & ~n3621;
  assign n3623 = n3622 ^ n2444;
  assign n3616 = n2634 ^ n2523;
  assign n3617 = n2524 & ~n3616;
  assign n3618 = n3617 ^ n2472;
  assign n3607 = ~n565 & ~n2371;
  assign n3608 = ~n2496 & ~n3607;
  assign n3609 = ~n2518 & ~n3608;
  assign n3610 = n3609 ^ n2350;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = n565 & n3611;
  assign n3613 = n3612 ^ n3610;
  assign n3600 = n573 & n2560;
  assign n3601 = n3600 ^ n2346;
  assign n3602 = n596 & ~n3601;
  assign n3603 = ~n2347 & ~n2488;
  assign n3604 = n2349 & n2492;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~n3602 & n3605;
  assign n3614 = n3613 ^ n3606;
  assign n3586 = n1108 & n2657;
  assign n3587 = n2344 & n2449;
  assign n3588 = ~n2345 & n2459;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3586 & n3589;
  assign n3591 = ~n595 & ~n3590;
  assign n3592 = n1108 & ~n2664;
  assign n3593 = n595 & n3589;
  assign n3594 = ~n3592 & n3593;
  assign n3595 = n1108 & n2656;
  assign n3596 = n2343 ^ n618;
  assign n3597 = n3595 & ~n3596;
  assign n3598 = ~n3594 & ~n3597;
  assign n3599 = ~n3591 & n3598;
  assign n3615 = n3614 ^ n3599;
  assign n3619 = n3618 ^ n3615;
  assign n3572 = n1451 & n2846;
  assign n3573 = ~n2360 & n2428;
  assign n3574 = n2342 & n2431;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = ~n3572 & n3575;
  assign n3577 = n812 & ~n3576;
  assign n3578 = n1451 & ~n2842;
  assign n3579 = ~n812 & n3575;
  assign n3580 = ~n3578 & n3579;
  assign n3581 = n1451 & n2841;
  assign n3582 = n2320 ^ n816;
  assign n3583 = n3581 & ~n3582;
  assign n3584 = ~n3580 & ~n3583;
  assign n3585 = ~n3577 & n3584;
  assign n3620 = n3619 ^ n3585;
  assign n3624 = n3623 ^ n3620;
  assign n3150 = n3095 ^ n3064;
  assign n3182 = ~n3128 & ~n3132;
  assign n3183 = n3182 ^ n2403;
  assign n3184 = ~n2384 & n3183;
  assign n3547 = n3150 & ~n3184;
  assign n3548 = n2845 & ~n3547;
  assign n3549 = ~n2407 & ~n2803;
  assign n3550 = n2318 & n2333;
  assign n3551 = n3550 ^ n30;
  assign n3552 = n3551 ^ n3550;
  assign n3553 = n2317 & n2329;
  assign n3554 = n3553 ^ n3550;
  assign n3555 = n3552 & n3554;
  assign n3556 = n3555 ^ n3550;
  assign n3557 = ~n3549 & ~n3556;
  assign n3558 = n3557 ^ n30;
  assign n3559 = ~n3548 & n3558;
  assign n3185 = n3184 ^ n3150;
  assign n3560 = ~n2795 & n3150;
  assign n3561 = n3560 ^ n30;
  assign n3562 = n2385 & n3561;
  assign n3563 = n3562 ^ n2938;
  assign n3564 = n3563 ^ n3562;
  assign n3565 = n3562 ^ n3184;
  assign n3566 = n3565 ^ n3562;
  assign n3567 = n3564 & n3566;
  assign n3568 = n3567 ^ n3562;
  assign n3569 = n3185 & n3568;
  assign n3570 = n3569 ^ n3562;
  assign n3571 = ~n3559 & ~n3570;
  assign n3625 = n3624 ^ n3571;
  assign n3629 = n3628 ^ n3625;
  assign n3667 = n3666 ^ n3629;
  assign n3144 = ~n3125 & ~n3143;
  assign n3145 = n3118 & ~n3144;
  assign n3146 = n3145 ^ x1;
  assign n3117 = n3116 ^ x22;
  assign n3147 = n3146 ^ n3117;
  assign n3098 = n3097 ^ n2321;
  assign n3099 = x1 & n3098;
  assign n3148 = n3147 ^ n3099;
  assign n3149 = n3148 ^ n3147;
  assign n3151 = n2322 & n3150;
  assign n3152 = n3151 ^ n3147;
  assign n3153 = n3152 ^ n3147;
  assign n3154 = ~n3149 & ~n3153;
  assign n3155 = n3154 ^ n3147;
  assign n3156 = ~x0 & ~n3155;
  assign n3157 = n3156 ^ n3147;
  assign n3045 = n3044 ^ n2420;
  assign n3158 = n3157 ^ n3045;
  assign n3159 = n3040 ^ n2823;
  assign n3161 = ~n3119 & ~n3126;
  assign n3162 = n3141 & ~n3161;
  assign n3163 = ~n3122 & ~n3162;
  assign n3164 = n3118 & n3163;
  assign n3165 = n3164 ^ n3097;
  assign n3160 = x1 & ~n3150;
  assign n3166 = n3165 ^ n3160;
  assign n3167 = n3166 ^ n3165;
  assign n3168 = n2322 & ~n2407;
  assign n3169 = n3168 ^ n3165;
  assign n3170 = n3169 ^ n3165;
  assign n3171 = ~n3167 & ~n3170;
  assign n3172 = n3171 ^ n3165;
  assign n3173 = ~x0 & n3172;
  assign n3174 = n3173 ^ n3165;
  assign n3175 = n3174 ^ n2327;
  assign n3496 = ~n3159 & n3175;
  assign n3539 = n3496 ^ n3045;
  assign n3540 = n3539 ^ n3045;
  assign n3177 = n3159 & ~n3175;
  assign n3218 = n2407 ^ n2327;
  assign n3217 = n2384 & n3118;
  assign n3219 = n3218 ^ n3217;
  assign n3215 = n2321 ^ n2317;
  assign n3216 = x1 & ~n3215;
  assign n3220 = n3219 ^ n3216;
  assign n3221 = n3220 ^ n3219;
  assign n3222 = n2320 & n2322;
  assign n3223 = n3222 ^ n3219;
  assign n3224 = n3223 ^ n3219;
  assign n3225 = ~n3221 & ~n3224;
  assign n3226 = n3225 ^ n3219;
  assign n3227 = ~x0 & n3226;
  assign n3228 = n3227 ^ n3219;
  assign n3214 = n3034 ^ n2881;
  assign n3229 = n3228 ^ n3214;
  assign n3243 = n3031 ^ n2897;
  assign n3231 = n2382 & n3118;
  assign n3232 = n3231 ^ n2317;
  assign n3230 = x1 & ~n2320;
  assign n3233 = n3232 ^ n3230;
  assign n3234 = n3233 ^ n3232;
  assign n3235 = n2322 & ~n2360;
  assign n3236 = n3235 ^ n3232;
  assign n3237 = n3236 ^ n3232;
  assign n3238 = ~n3234 & ~n3237;
  assign n3239 = n3238 ^ n3232;
  assign n3240 = ~x0 & ~n3239;
  assign n3241 = n3240 ^ n3232;
  assign n3242 = n3241 ^ n2327;
  assign n3244 = n3243 ^ n3242;
  assign n3254 = n3028 ^ n2919;
  assign n3245 = n2841 & n3118;
  assign n3246 = n3245 ^ n2320;
  assign n3247 = x0 & ~n3246;
  assign n3248 = ~n2360 & n3188;
  assign n3250 = n2342 & n3249;
  assign n3251 = ~n3248 & ~n3250;
  assign n3252 = ~n3247 & n3251;
  assign n3253 = n3252 ^ n2327;
  assign n3255 = n3254 ^ n3253;
  assign n3256 = n3022 ^ n2970;
  assign n3265 = n3019 ^ n3009;
  assign n3257 = n2656 & n3118;
  assign n3258 = n3257 ^ n2343;
  assign n3259 = x0 & ~n3258;
  assign n3260 = n2344 & n3188;
  assign n3261 = ~n2345 & n3249;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = ~n3259 & n3262;
  assign n3264 = n3263 ^ n2327;
  assign n3266 = n3265 ^ n3264;
  assign n3285 = n30 & ~n2995;
  assign n3286 = n3285 ^ n2977;
  assign n3283 = n2977 & ~n2995;
  assign n3284 = n3283 ^ n1100;
  assign n3287 = n3286 ^ n3284;
  assign n3288 = n2371 & n3287;
  assign n3289 = n3288 ^ n3284;
  assign n3268 = n2344 & n3267;
  assign n3269 = ~n2345 & n3188;
  assign n3270 = ~n2346 & n3249;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = ~n3268 & n3271;
  assign n3273 = n2327 & n3272;
  assign n3274 = n2445 ^ n2344;
  assign n3275 = n3206 & n3274;
  assign n3276 = n3273 & ~n3275;
  assign n3277 = n2323 & ~n3272;
  assign n3278 = n2322 & n2325;
  assign n3279 = ~n3181 & ~n3278;
  assign n3280 = n3274 & ~n3279;
  assign n3281 = ~n3277 & ~n3280;
  assign n3282 = ~n3276 & n3281;
  assign n3290 = n3289 ^ n3282;
  assign n3317 = n2864 ^ n32;
  assign n3318 = n3317 ^ n2327;
  assign n3319 = n2865 ^ n2327;
  assign n3320 = n2350 ^ n2327;
  assign n3321 = n3320 ^ n2327;
  assign n3322 = n3319 & n3321;
  assign n3323 = n3322 ^ n2327;
  assign n3324 = n3318 & ~n3323;
  assign n3325 = n3324 ^ n2864;
  assign n3291 = n2350 & n2385;
  assign n3326 = n3325 ^ n3291;
  assign n3327 = n3291 ^ n32;
  assign n3328 = n3291 ^ n2371;
  assign n3329 = n3291 & ~n3328;
  assign n3330 = n3329 ^ n3291;
  assign n3331 = ~n3327 & n3330;
  assign n3332 = n3331 ^ n3329;
  assign n3333 = n3332 ^ n3291;
  assign n3334 = n3333 ^ n2371;
  assign n3335 = n3326 & ~n3334;
  assign n3336 = n3335 ^ n3291;
  assign n3296 = n2500 & n3118;
  assign n3297 = n3296 ^ n2347;
  assign n3298 = x0 & ~n3297;
  assign n3299 = n2349 & n3188;
  assign n3300 = n2350 & n3249;
  assign n3301 = ~n3299 & ~n3300;
  assign n3302 = ~n3298 & n3301;
  assign n3312 = n1323 & ~n2327;
  assign n3313 = ~n2371 & n3312;
  assign n3303 = n2349 ^ n1323;
  assign n3304 = n3303 ^ n1323;
  assign n3305 = n2204 ^ n1323;
  assign n3306 = n3305 ^ n1323;
  assign n3307 = ~n3304 & ~n3306;
  assign n3308 = n3307 ^ n1323;
  assign n3309 = n2371 & ~n3308;
  assign n3310 = n3309 ^ n1323;
  assign n3311 = n2327 & ~n3310;
  assign n3314 = n3313 ^ n3311;
  assign n3315 = ~n3302 & n3314;
  assign n3316 = n3315 ^ n3311;
  assign n3337 = n3336 ^ n3316;
  assign n3338 = x0 & n2346;
  assign n3339 = n2347 & n3188;
  assign n3340 = n2322 & ~n2349;
  assign n3341 = x0 & n3118;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = ~n3339 & n3342;
  assign n3344 = ~n3338 & n3343;
  assign n3345 = n2324 & ~n3344;
  assign n3207 = n3206 ^ n2326;
  assign n3346 = ~n2743 & n3207;
  assign n3347 = n3346 ^ n2326;
  assign n3348 = n3345 & ~n3347;
  assign n3187 = ~n25 & n2323;
  assign n3349 = n3187 & n3344;
  assign n3350 = ~n2743 & n3181;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n3348 & n3351;
  assign n3353 = n3352 ^ n3336;
  assign n3354 = n3337 & n3353;
  assign n3355 = n3354 ^ n3316;
  assign n3292 = n2371 & ~n3291;
  assign n3293 = n30 & ~n2866;
  assign n3294 = ~n3292 & n3293;
  assign n3295 = n3294 ^ n2994;
  assign n3356 = n3355 ^ n3295;
  assign n3357 = ~n2345 & n3267;
  assign n3358 = ~n2346 & n3188;
  assign n3359 = ~n2347 & n3249;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~n3357 & n3360;
  assign n3362 = n2327 & n3361;
  assign n3363 = n2525 ^ n2345;
  assign n3364 = n3341 & ~n3363;
  assign n3365 = n3362 & ~n3364;
  assign n3366 = n2323 & ~n3361;
  assign n3367 = ~n3279 & ~n3363;
  assign n3368 = ~n3366 & ~n3367;
  assign n3369 = ~n3365 & n3368;
  assign n3370 = n3369 ^ n3295;
  assign n3371 = n3356 & n3370;
  assign n3372 = n3371 ^ n3355;
  assign n3373 = n3372 ^ n3289;
  assign n3374 = n3290 & n3373;
  assign n3375 = n3374 ^ n3282;
  assign n3376 = n3375 ^ n3265;
  assign n3377 = n3266 & ~n3376;
  assign n3378 = n3377 ^ n3264;
  assign n3379 = n3256 & ~n3378;
  assign n3382 = n2322 & n2344;
  assign n3380 = n2637 & n3118;
  assign n3381 = n3380 ^ n2342;
  assign n3383 = n3382 ^ n3381;
  assign n3384 = n3383 ^ n3381;
  assign n3385 = x1 & ~n2343;
  assign n3386 = n3385 ^ n3381;
  assign n3387 = n3386 ^ n3381;
  assign n3388 = ~n3384 & ~n3387;
  assign n3389 = n3388 ^ n3381;
  assign n3390 = ~x0 & ~n3389;
  assign n3391 = n3390 ^ n3381;
  assign n3392 = n3391 ^ n2327;
  assign n3393 = n3025 ^ n2953;
  assign n3394 = n2421 & n3118;
  assign n3395 = n3394 ^ n2360;
  assign n3396 = x0 & ~n3395;
  assign n3397 = n2342 & n3188;
  assign n3398 = ~n2343 & n3249;
  assign n3399 = ~n3397 & ~n3398;
  assign n3400 = ~n3396 & n3399;
  assign n3401 = n3400 ^ n3391;
  assign n3402 = ~n3393 & ~n3401;
  assign n3403 = ~n3392 & n3402;
  assign n3404 = n3403 ^ n3392;
  assign n3405 = ~n3379 & ~n3404;
  assign n3406 = n3400 ^ n2327;
  assign n3407 = n3406 ^ n3393;
  assign n3408 = ~n3256 & n3378;
  assign n3409 = n3408 ^ n3406;
  assign n3410 = n3407 & ~n3409;
  assign n3411 = n3410 ^ n3393;
  assign n3412 = ~n3405 & ~n3411;
  assign n3413 = n3412 ^ n3254;
  assign n3414 = ~n3255 & ~n3413;
  assign n3415 = n3414 ^ n3253;
  assign n3416 = n3415 ^ n3243;
  assign n3417 = n3244 & n3416;
  assign n3418 = n3417 ^ n3242;
  assign n3419 = n3418 ^ n3214;
  assign n3420 = n3229 & n3419;
  assign n3421 = n3420 ^ n3228;
  assign n3186 = n3181 & ~n3185;
  assign n3189 = ~n3118 & ~n3188;
  assign n3190 = ~n3150 & n3189;
  assign n3191 = ~n2317 & n2322;
  assign n3192 = x1 ^ x0;
  assign n3193 = x1 & ~n3192;
  assign n3194 = n3193 ^ x1;
  assign n3195 = n2407 ^ x1;
  assign n3196 = n3194 & n3195;
  assign n3197 = n3196 ^ n3193;
  assign n3198 = n3197 ^ x1;
  assign n3199 = n3198 ^ x0;
  assign n3200 = ~n3191 & ~n3199;
  assign n3201 = ~n3190 & ~n3200;
  assign n3202 = n3187 & ~n3201;
  assign n3203 = ~n3186 & ~n3202;
  assign n3204 = n2324 & n3201;
  assign n3208 = n3206 ^ n3185;
  assign n3209 = n3208 ^ n3206;
  assign n3210 = n3207 & n3209;
  assign n3211 = n3210 ^ n3206;
  assign n3212 = n3204 & ~n3211;
  assign n3213 = n3203 & ~n3212;
  assign n3422 = n3421 ^ n3213;
  assign n3423 = n3037 ^ n2861;
  assign n3424 = n3423 ^ n3213;
  assign n3425 = n3422 & ~n3424;
  assign n3426 = n3425 ^ n3421;
  assign n3499 = ~n3177 & n3426;
  assign n3541 = n3499 ^ n3045;
  assign n3542 = n3541 ^ n3045;
  assign n3543 = ~n3540 & ~n3542;
  assign n3544 = n3543 ^ n3045;
  assign n3545 = n3158 & ~n3544;
  assign n3546 = n3545 ^ n3157;
  assign n3782 = n3666 ^ n3546;
  assign n3783 = ~n3667 & ~n3782;
  assign n3784 = n3783 ^ n3546;
  assign n3760 = n2795 & n3163;
  assign n3761 = n3760 ^ n30;
  assign n3762 = n3761 ^ n3097;
  assign n3763 = n2385 & n3762;
  assign n3764 = n2329 ^ n30;
  assign n3765 = n2407 ^ n2329;
  assign n3766 = n2329 & n3765;
  assign n3767 = n3766 ^ n2329;
  assign n3768 = ~n3764 & n3767;
  assign n3769 = n3768 ^ n3766;
  assign n3770 = n3769 ^ n2329;
  assign n3771 = n3770 ^ n2407;
  assign n3772 = n2808 & n3771;
  assign n3773 = n3772 ^ n2329;
  assign n3774 = n3150 ^ n2801;
  assign n3775 = n3774 ^ n2801;
  assign n3776 = n2805 & ~n3775;
  assign n3777 = n3776 ^ n2801;
  assign n3778 = ~n3773 & ~n3777;
  assign n3779 = ~n3763 & n3778;
  assign n3756 = n3628 ^ n3571;
  assign n3757 = n3625 & n3756;
  assign n3758 = n3757 ^ n3628;
  assign n3751 = n3623 ^ n3585;
  assign n3752 = n3620 & n3751;
  assign n3753 = n3752 ^ n3623;
  assign n3747 = n3618 ^ n3614;
  assign n3748 = ~n3615 & ~n3747;
  assign n3749 = n3748 ^ n3599;
  assign n3738 = n573 & n2525;
  assign n3739 = n3738 ^ n2345;
  assign n3740 = n596 & ~n3739;
  assign n3741 = ~n2346 & ~n2488;
  assign n3742 = ~n2347 & n2492;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = ~n3740 & n3743;
  assign n3733 = n3609 ^ n3606;
  assign n3734 = n3610 & ~n3733;
  assign n3735 = n3734 ^ n2350;
  assign n3736 = n3735 ^ n2349;
  assign n3737 = ~n565 & ~n3736;
  assign n3745 = n3744 ^ n3737;
  assign n3719 = n1108 & n2638;
  assign n3720 = ~n2343 & n2449;
  assign n3721 = n2344 & n2459;
  assign n3722 = ~n3720 & ~n3721;
  assign n3723 = ~n3719 & n3722;
  assign n3724 = ~n595 & ~n3723;
  assign n3725 = n1108 & ~n2645;
  assign n3726 = n595 & n3722;
  assign n3727 = ~n3725 & n3726;
  assign n3728 = n1108 & n2637;
  assign n3729 = n2342 ^ n618;
  assign n3730 = n3728 & n3729;
  assign n3731 = ~n3727 & ~n3730;
  assign n3732 = ~n3724 & n3731;
  assign n3746 = n3745 ^ n3732;
  assign n3750 = n3749 ^ n3746;
  assign n3754 = n3753 ^ n3750;
  assign n3703 = n2317 & ~n2382;
  assign n3704 = n1451 & n3703;
  assign n3705 = ~n2320 & n2428;
  assign n3706 = ~n2360 & n2431;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = ~n3704 & n3707;
  assign n3709 = n812 & ~n3708;
  assign n3710 = ~n2317 & ~n2382;
  assign n3711 = n1451 & ~n3710;
  assign n3712 = ~n812 & n3707;
  assign n3713 = ~n3711 & n3712;
  assign n3714 = n1451 & n2382;
  assign n3715 = n2317 ^ n816;
  assign n3716 = n3714 & n3715;
  assign n3717 = ~n3713 & ~n3716;
  assign n3718 = ~n3709 & n3717;
  assign n3755 = n3754 ^ n3718;
  assign n3759 = n3758 ^ n3755;
  assign n3780 = n3779 ^ n3759;
  assign n3678 = n124 & n638;
  assign n3679 = n60 & ~n3678;
  assign n3680 = ~n326 & ~n459;
  assign n3681 = n94 & ~n136;
  assign n3682 = n3680 & ~n3681;
  assign n3683 = ~n3679 & n3682;
  assign n3684 = ~n199 & ~n676;
  assign n3685 = n3683 & n3684;
  assign n3686 = ~n228 & ~n367;
  assign n3687 = n342 & n3686;
  assign n3688 = n94 & ~n3637;
  assign n3689 = n3687 & ~n3688;
  assign n3690 = n3685 & n3689;
  assign n3691 = n1082 & n3690;
  assign n3674 = n3642 & n3654;
  assign n3675 = n3643 & ~n3651;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = n3118 & n3676;
  assign n3692 = n3691 ^ n3677;
  assign n3673 = x1 & n3643;
  assign n3693 = n3692 ^ n3673;
  assign n3694 = n3693 ^ n3692;
  assign n3695 = n2322 & ~n3116;
  assign n3696 = n3695 ^ n3692;
  assign n3697 = n3696 ^ n3692;
  assign n3698 = ~n3694 & ~n3697;
  assign n3699 = n3698 ^ n3692;
  assign n3700 = ~x0 & n3699;
  assign n3701 = n3700 ^ n3692;
  assign n3702 = n3701 ^ n2327;
  assign n3781 = n3780 ^ n3702;
  assign n3785 = n3784 ^ n3781;
  assign n3795 = n3794 ^ n3785;
  assign n3176 = n3175 ^ n3159;
  assign n3178 = n3177 ^ n3176;
  assign n3427 = ~n445 & ~n845;
  assign n3428 = ~n397 & n3427;
  assign n3429 = n2279 & n3428;
  assign n3430 = n2038 & n3429;
  assign n3431 = ~n416 & ~n1043;
  assign n3432 = n3430 & n3431;
  assign n3433 = ~n414 & n3432;
  assign n3434 = ~n180 & ~n214;
  assign n3435 = ~n111 & n3434;
  assign n3436 = n171 & ~n336;
  assign n3437 = n2115 & ~n3436;
  assign n3438 = n3435 & n3437;
  assign n3439 = n2125 & n3438;
  assign n3440 = n250 & ~n681;
  assign n3441 = n2232 & n3440;
  assign n3442 = n3439 & n3441;
  assign n3443 = n172 & ~n349;
  assign n3444 = n273 & ~n3443;
  assign n3445 = n645 & n3444;
  assign n3446 = n3442 & n3445;
  assign n3447 = n3433 & n3446;
  assign n3448 = ~n3426 & ~n3447;
  assign n3449 = ~n60 & ~n438;
  assign n3450 = ~n187 & n3449;
  assign n3451 = n178 & n351;
  assign n3452 = ~n3450 & ~n3451;
  assign n3453 = n1060 & ~n3452;
  assign n3456 = ~n327 & ~n676;
  assign n3457 = n3455 & n3456;
  assign n3458 = n182 & n3457;
  assign n3459 = n3453 & n3458;
  assign n3460 = ~n215 & ~n622;
  assign n3461 = n658 & n3460;
  assign n3462 = n3459 & n3461;
  assign n3463 = ~n107 & ~n436;
  assign n3464 = n3079 & n3463;
  assign n3465 = n927 & n3464;
  assign n3466 = ~n95 & n166;
  assign n3467 = ~n106 & n3466;
  assign n3468 = ~n629 & ~n3467;
  assign n3469 = ~n709 & ~n3468;
  assign n3470 = n3465 & n3469;
  assign n3471 = n2176 & n3470;
  assign n3472 = ~n111 & ~n186;
  assign n3473 = n60 & ~n349;
  assign n3474 = ~n727 & ~n3473;
  assign n3475 = n3472 & n3474;
  assign n3476 = n493 & n2237;
  assign n3477 = n3475 & n3476;
  assign n3478 = ~n464 & ~n647;
  assign n3479 = n184 & ~n309;
  assign n3480 = ~n1964 & ~n3479;
  assign n3481 = n3478 & n3480;
  assign n3482 = n3477 & n3481;
  assign n3483 = n3471 & n3482;
  assign n3484 = n3462 & n3483;
  assign n3485 = n3448 & ~n3484;
  assign n3486 = n3485 ^ n3176;
  assign n3487 = n3486 ^ n3485;
  assign n3488 = n3485 ^ n3426;
  assign n3489 = ~n3487 & ~n3488;
  assign n3490 = n3489 ^ n3485;
  assign n3491 = ~n3178 & n3490;
  assign n3492 = n3491 ^ n3177;
  assign n3493 = n3158 & ~n3492;
  assign n3494 = ~n3177 & n3484;
  assign n3495 = ~n3158 & ~n3494;
  assign n3497 = ~n3448 & n3496;
  assign n3498 = n3495 & ~n3497;
  assign n3500 = n3447 & n3499;
  assign n3501 = n3498 & ~n3500;
  assign n3502 = ~n3493 & ~n3501;
  assign n3503 = ~n3176 & ~n3447;
  assign n3504 = ~n3448 & n3484;
  assign n3505 = ~n3503 & n3504;
  assign n3506 = ~n3502 & ~n3505;
  assign n3507 = ~n163 & ~n2030;
  assign n3508 = ~n659 & ~n2123;
  assign n3509 = ~n298 & ~n398;
  assign n3510 = n3508 & n3509;
  assign n3511 = n900 & n3510;
  assign n3512 = n2036 & n3059;
  assign n3513 = n184 & ~n2389;
  assign n3514 = ~n443 & ~n3513;
  assign n3515 = ~n71 & n171;
  assign n3516 = ~n721 & ~n3515;
  assign n3517 = ~n314 & n3516;
  assign n3518 = n3514 & n3517;
  assign n3519 = n3512 & n3518;
  assign n3520 = n3511 & n3519;
  assign n3521 = n671 & n3520;
  assign n3522 = ~n3507 & n3521;
  assign n3523 = n487 & ~n539;
  assign n3524 = ~n355 & ~n491;
  assign n3525 = n60 & ~n115;
  assign n3526 = ~n654 & ~n3525;
  assign n3527 = n3524 & n3526;
  assign n3528 = n3091 & n3527;
  assign n3529 = n530 & n3528;
  assign n3530 = n276 & n3068;
  assign n3531 = ~n227 & n634;
  assign n3532 = n437 & n3531;
  assign n3533 = n1973 & n3532;
  assign n3534 = n3530 & n3533;
  assign n3535 = n3529 & n3534;
  assign n3536 = n3523 & n3535;
  assign n3537 = n3522 & n3536;
  assign n3538 = n3506 & ~n3537;
  assign n3668 = n3667 ^ n3546;
  assign n3669 = n3538 & n3668;
  assign n3670 = ~n3506 & n3537;
  assign n3671 = ~n3668 & n3670;
  assign n3672 = ~n3669 & ~n3671;
  assign n3796 = n3795 ^ n3672;
  assign n3948 = ~n465 & ~n676;
  assign n3949 = n172 & ~n422;
  assign n3950 = ~n375 & ~n3949;
  assign n3951 = n3948 & n3950;
  assign n3952 = n3068 & n3951;
  assign n3953 = n60 & ~n3085;
  assign n3954 = ~n278 & ~n3953;
  assign n3955 = n3427 & n3954;
  assign n3956 = n3952 & n3955;
  assign n3957 = n2019 & n3956;
  assign n3958 = n415 & ~n674;
  assign n3959 = ~n107 & ~n399;
  assign n3960 = n3958 & n3959;
  assign n3961 = n3957 & n3960;
  assign n3962 = n3520 & n3961;
  assign n3817 = ~n628 & ~n887;
  assign n3818 = ~n214 & n3817;
  assign n3963 = n3106 & n3818;
  assign n3964 = n3530 & n3963;
  assign n3965 = ~n708 & ~n3964;
  assign n3966 = ~n131 & ~n1012;
  assign n3967 = ~n3965 & n3966;
  assign n3968 = n3962 & n3967;
  assign n3944 = n3784 ^ n3702;
  assign n3945 = ~n3781 & ~n3944;
  assign n3946 = n3945 ^ n3784;
  assign n3939 = n3779 ^ n3755;
  assign n3940 = ~n3759 & n3939;
  assign n3941 = n3940 ^ n3758;
  assign n3934 = n3753 ^ n3718;
  assign n3935 = n3754 & n3934;
  assign n3936 = n3935 ^ n3718;
  assign n3929 = n3749 ^ n3745;
  assign n3930 = n3746 & ~n3929;
  assign n3931 = n3930 ^ n3732;
  assign n3903 = n572 & ~n2345;
  assign n3904 = n3903 ^ n579;
  assign n3905 = n3904 ^ n3903;
  assign n3906 = ~n2346 & n2504;
  assign n3907 = n3906 ^ n3903;
  assign n3908 = ~n3905 & n3907;
  assign n3909 = n3908 ^ n3903;
  assign n3901 = n573 & n2445;
  assign n3902 = n3901 ^ n2344;
  assign n3910 = n3909 ^ n3902;
  assign n3911 = n3910 ^ n3902;
  assign n3912 = n2346 ^ n2345;
  assign n3913 = n3912 ^ n2345;
  assign n3914 = n2345 ^ n565;
  assign n3915 = n3914 ^ n2345;
  assign n3916 = ~n3913 & n3915;
  assign n3917 = n3916 ^ n2345;
  assign n3918 = n595 & ~n3917;
  assign n3919 = n3918 ^ n2345;
  assign n3920 = ~n572 & ~n3919;
  assign n3921 = n3920 ^ n3902;
  assign n3922 = n3921 ^ n3902;
  assign n3923 = ~n3911 & ~n3922;
  assign n3924 = n3923 ^ n3902;
  assign n3925 = ~n596 & ~n3924;
  assign n3926 = n3925 ^ n3902;
  assign n3895 = n3744 ^ n2349;
  assign n3896 = n3736 & n3895;
  assign n3897 = n3896 ^ n2349;
  assign n3898 = ~n565 & n3897;
  assign n3899 = n3898 ^ n2347;
  assign n3900 = ~n565 & n3899;
  assign n3927 = n3926 ^ n3900;
  assign n3875 = n2360 ^ n618;
  assign n3876 = n1108 & n2421;
  assign n3877 = n3875 & n3876;
  assign n3878 = n2342 & n2449;
  assign n3879 = ~n2343 & n2459;
  assign n3880 = ~n3878 & ~n3879;
  assign n3881 = n3880 ^ n595;
  assign n3882 = n1108 & ~n2436;
  assign n3883 = n3882 ^ n3880;
  assign n3884 = n2422 & n2464;
  assign n3885 = n3884 ^ n3882;
  assign n3886 = n3882 & ~n3885;
  assign n3887 = n3886 ^ n3882;
  assign n3888 = n3883 & n3887;
  assign n3889 = n3888 ^ n3886;
  assign n3890 = n3889 ^ n3882;
  assign n3891 = n3890 ^ n3884;
  assign n3892 = n3881 & ~n3891;
  assign n3893 = n3892 ^ n3884;
  assign n3894 = ~n3877 & ~n3893;
  assign n3928 = n3927 ^ n3894;
  assign n3932 = n3931 ^ n3928;
  assign n3861 = n1451 & n2413;
  assign n3862 = n2317 & n2428;
  assign n3863 = ~n2320 & n2431;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = ~n3861 & n3864;
  assign n3866 = ~n812 & ~n3865;
  assign n3867 = n1451 & ~n2417;
  assign n3868 = n812 & n3864;
  assign n3869 = ~n3867 & n3868;
  assign n3870 = n2407 ^ n816;
  assign n3871 = n1451 & n3870;
  assign n3872 = n2384 & n3871;
  assign n3873 = ~n3869 & ~n3872;
  assign n3874 = ~n3866 & n3873;
  assign n3933 = n3932 ^ n3874;
  assign n3937 = n3936 ^ n3933;
  assign n3845 = ~n3116 & ~n3144;
  assign n3846 = n2412 & n3845;
  assign n3847 = ~n2803 & ~n3097;
  assign n3848 = n2867 & ~n3150;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n30 & ~n3849;
  assign n3851 = ~n3846 & ~n3850;
  assign n3852 = n2385 & n3144;
  assign n3853 = n3116 ^ n32;
  assign n3854 = n3852 & n3853;
  assign n3855 = n3851 & ~n3854;
  assign n3856 = n3116 & ~n3144;
  assign n3857 = n2385 & ~n3856;
  assign n3858 = ~n30 & n3849;
  assign n3859 = ~n3857 & n3858;
  assign n3860 = n3855 & ~n3859;
  assign n3938 = n3937 ^ n3860;
  assign n3942 = n3941 ^ n3938;
  assign n3819 = n95 & ~n1057;
  assign n3820 = n3818 & ~n3819;
  assign n3821 = n1299 & n3820;
  assign n3822 = n328 & n2076;
  assign n3823 = n3821 & n3822;
  assign n3824 = n304 & n626;
  assign n3825 = n106 & ~n3824;
  assign n3826 = n543 & ~n3825;
  assign n3827 = ~n102 & n2283;
  assign n3828 = ~n654 & n3827;
  assign n3829 = ~n674 & n3828;
  assign n3830 = n3826 & n3829;
  assign n3831 = n646 & n3830;
  assign n3832 = n3823 & n3831;
  assign n3833 = n2254 & n3832;
  assign n3813 = ~n3674 & ~n3691;
  assign n3814 = ~n3675 & n3691;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3118 & n3815;
  assign n3834 = n3833 ^ n3816;
  assign n3812 = n2322 & n3643;
  assign n3835 = n3834 ^ n3812;
  assign n3836 = n3835 ^ n3834;
  assign n3837 = x1 & ~n3691;
  assign n3838 = n3837 ^ n3834;
  assign n3839 = n3838 ^ n3834;
  assign n3840 = ~n3836 & ~n3839;
  assign n3841 = n3840 ^ n3834;
  assign n3842 = ~x0 & n3841;
  assign n3843 = n3842 ^ n3834;
  assign n3844 = n3843 ^ n2327;
  assign n3943 = n3942 ^ n3844;
  assign n3947 = n3946 ^ n3943;
  assign n3969 = n3968 ^ n3947;
  assign n3797 = x23 ^ x22;
  assign n3798 = n3797 ^ n3794;
  assign n3799 = ~n3795 & n3798;
  assign n3800 = n3799 ^ n3785;
  assign n3801 = n3671 & ~n3800;
  assign n3802 = ~n3785 & n3794;
  assign n3803 = ~n3797 & n3802;
  assign n3804 = n3803 ^ n3800;
  assign n3805 = ~n3669 & n3804;
  assign n3806 = n3805 ^ n3800;
  assign n3807 = ~n3801 & ~n3806;
  assign n3808 = n3785 & ~n3794;
  assign n3809 = ~n3671 & n3808;
  assign n3810 = n3797 & n3809;
  assign n3811 = n3807 & ~n3810;
  assign n3970 = n3969 ^ n3811;
  assign n3988 = ~n3802 & n3969;
  assign n3989 = n3669 & ~n3988;
  assign n3971 = n3537 ^ n3506;
  assign n3972 = n3668 ^ n3537;
  assign n3973 = ~n3971 & n3972;
  assign n3974 = n3973 ^ n3506;
  assign n3990 = ~n3671 & ~n3795;
  assign n3991 = ~n3974 & n3990;
  assign n3992 = ~n3989 & ~n3991;
  assign n3993 = n3669 & n3808;
  assign n3994 = ~n3969 & ~n3993;
  assign n3995 = ~n3992 & ~n3994;
  assign n3975 = ~n3802 & n3974;
  assign n3976 = ~n3669 & n3975;
  assign n3977 = ~n3808 & n3969;
  assign n3978 = ~n3976 & n3977;
  assign n3979 = n3969 ^ n3671;
  assign n3980 = n3808 ^ n3802;
  assign n3981 = n3969 ^ n3808;
  assign n3982 = n3981 ^ n3808;
  assign n3983 = n3980 & ~n3982;
  assign n3984 = n3983 ^ n3808;
  assign n3985 = n3979 & ~n3984;
  assign n3986 = n3985 ^ n3671;
  assign n3987 = ~n3978 & n3986;
  assign n3996 = n3995 ^ n3987;
  assign n4151 = n3946 ^ n3844;
  assign n4152 = n3943 & ~n4151;
  assign n4153 = n4152 ^ n3946;
  assign n4146 = n3941 ^ n3860;
  assign n4147 = ~n3938 & n4146;
  assign n4148 = n4147 ^ n3941;
  assign n4142 = n3936 ^ n3932;
  assign n4143 = n3933 & n4142;
  assign n4144 = n4143 ^ n3874;
  assign n4137 = n3931 ^ n3927;
  assign n4138 = n3928 & n4137;
  assign n4139 = n4138 ^ n3894;
  assign n4128 = n573 & n2656;
  assign n4129 = n4128 ^ n2343;
  assign n4130 = n596 & ~n4129;
  assign n4131 = n2344 & ~n2488;
  assign n4132 = ~n2345 & n2492;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = ~n4130 & n4133;
  assign n4123 = n3926 ^ n3898;
  assign n4124 = ~n3899 & n4123;
  assign n4125 = n4124 ^ n2347;
  assign n4126 = n4125 ^ n2346;
  assign n4127 = ~n565 & ~n4126;
  assign n4135 = n4134 ^ n4127;
  assign n4109 = n2320 ^ n618;
  assign n4110 = n1108 & n2841;
  assign n4111 = n4109 & n4110;
  assign n4112 = ~n2360 & n2449;
  assign n4113 = n2342 & n2459;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = n4114 ^ n595;
  assign n4117 = n1108 & ~n2842;
  assign n4118 = ~n595 & n4117;
  assign n4116 = n2464 & n2846;
  assign n4119 = n4118 ^ n4116;
  assign n4120 = n4115 & ~n4119;
  assign n4121 = n4120 ^ n4116;
  assign n4122 = ~n4111 & ~n4121;
  assign n4136 = n4135 ^ n4122;
  assign n4140 = n4139 ^ n4136;
  assign n4082 = n2407 ^ n812;
  assign n4083 = n2425 & ~n4082;
  assign n4084 = n2317 ^ n812;
  assign n4085 = ~n812 & n817;
  assign n4086 = n4085 ^ n812;
  assign n4087 = n4084 & ~n4086;
  assign n4088 = n4087 ^ n4085;
  assign n4089 = n4088 ^ n812;
  assign n4090 = n4089 ^ n816;
  assign n4091 = n2424 & n4090;
  assign n4092 = n4091 ^ n816;
  assign n4093 = ~n4083 & ~n4092;
  assign n4094 = ~n812 & n2424;
  assign n4095 = ~n2407 & n4094;
  assign n4096 = n812 & n2425;
  assign n4097 = ~n2317 & n4096;
  assign n4098 = n816 & ~n4097;
  assign n4099 = ~n4095 & n4098;
  assign n4100 = ~n4093 & ~n4099;
  assign n4101 = n812 & n2407;
  assign n4102 = n2424 & n4101;
  assign n4103 = ~n4100 & ~n4102;
  assign n4104 = ~n817 & n3184;
  assign n4105 = n4104 ^ n812;
  assign n4106 = n4105 ^ n3150;
  assign n4107 = n1451 & ~n4106;
  assign n4108 = n4103 & ~n4107;
  assign n4141 = n4140 ^ n4108;
  assign n4145 = n4144 ^ n4141;
  assign n4149 = n4148 ^ n4145;
  assign n4064 = n3814 ^ n3813;
  assign n4065 = ~n3833 & n4064;
  assign n4066 = n4065 ^ n3813;
  assign n4067 = n4066 ^ n3205;
  assign n4068 = n4067 ^ n3205;
  assign n4069 = n3205 ^ n2321;
  assign n4070 = ~n4068 & n4069;
  assign n4071 = n4070 ^ n3205;
  assign n4062 = n3833 ^ n2321;
  assign n4063 = x1 & n4062;
  assign n4072 = n4071 ^ n4063;
  assign n4073 = n4072 ^ n4071;
  assign n4074 = n2322 & n3691;
  assign n4075 = n4074 ^ n4071;
  assign n4076 = n4075 ^ n4071;
  assign n4077 = ~n4073 & ~n4076;
  assign n4078 = n4077 ^ n4071;
  assign n4079 = ~x0 & n4078;
  assign n4080 = n4079 ^ n4071;
  assign n4022 = n32 & n3655;
  assign n4023 = n3643 & ~n4022;
  assign n4024 = n3116 ^ n30;
  assign n4025 = n4024 ^ n3116;
  assign n4026 = n3116 ^ n3097;
  assign n4027 = n4026 ^ n3116;
  assign n4028 = n4025 & ~n4027;
  assign n4029 = n4028 ^ n3116;
  assign n4030 = ~n32 & ~n4029;
  assign n4031 = n4030 ^ n3116;
  assign n4032 = n2328 & ~n4031;
  assign n4033 = n2334 & ~n3116;
  assign n4034 = n2337 & ~n3097;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = ~n4032 & n4035;
  assign n4037 = n4036 ^ n2385;
  assign n4038 = n4037 ^ n2385;
  assign n4039 = n3655 ^ n2385;
  assign n4040 = n4039 ^ n2385;
  assign n4041 = n4038 & n4040;
  assign n4042 = n4041 ^ n2385;
  assign n4043 = n30 & n4042;
  assign n4044 = n4043 ^ n2385;
  assign n4045 = n4023 & n4044;
  assign n4046 = n4036 ^ n30;
  assign n4047 = ~n3643 & ~n3655;
  assign n4048 = n2385 & ~n4047;
  assign n4049 = n4048 ^ n30;
  assign n4050 = ~n3643 & n3655;
  assign n4051 = n2938 & n4050;
  assign n4052 = n4051 ^ n30;
  assign n4053 = n30 & ~n4052;
  assign n4054 = n4053 ^ n30;
  assign n4055 = n4049 & n4054;
  assign n4056 = n4055 ^ n4053;
  assign n4057 = n4056 ^ n30;
  assign n4058 = n4057 ^ n4051;
  assign n4059 = ~n4046 & ~n4058;
  assign n4060 = n4059 ^ n4051;
  assign n4061 = ~n4045 & ~n4060;
  assign n4081 = n4080 ^ n4061;
  assign n4150 = n4149 ^ n4081;
  assign n4154 = n4153 ^ n4150;
  assign n4155 = n4154 ^ n3995;
  assign n4005 = n101 & n349;
  assign n4006 = n106 & ~n4005;
  assign n4007 = ~n1964 & ~n4006;
  assign n4008 = ~n232 & ~n444;
  assign n4009 = n4007 & n4008;
  assign n4010 = ~n255 & ~n278;
  assign n4011 = n370 & n4010;
  assign n4012 = n4009 & n4011;
  assign n4013 = ~n434 & ~n479;
  assign n4014 = n159 & n838;
  assign n4015 = n110 & ~n4014;
  assign n4016 = ~n260 & ~n398;
  assign n4017 = ~n4015 & n4016;
  assign n4018 = n4013 & n4017;
  assign n4019 = n4012 & n4018;
  assign n4020 = n637 & n4019;
  assign n4021 = n3433 & n4020;
  assign n4156 = n4155 ^ n4021;
  assign n3997 = n3975 ^ n3968;
  assign n3998 = n3997 ^ n3968;
  assign n3999 = n3968 ^ n3808;
  assign n4000 = n3999 ^ n3968;
  assign n4001 = ~n3998 & ~n4000;
  assign n4002 = n4001 ^ n3968;
  assign n4003 = n3969 & ~n4002;
  assign n4004 = n4003 ^ n3947;
  assign n4157 = n4156 ^ n4004;
  assign n4158 = n4157 ^ n3987;
  assign n4159 = n4158 ^ n4157;
  assign n4160 = n4157 ^ n3797;
  assign n4161 = ~n4159 & n4160;
  assign n4162 = n4161 ^ n4157;
  assign n4163 = ~n3996 & n4162;
  assign n4164 = n4163 ^ n4157;
  assign n4336 = n2079 & n3959;
  assign n4337 = ~n235 & ~n326;
  assign n4338 = n4336 & n4337;
  assign n4339 = ~n180 & ~n264;
  assign n4340 = ~n229 & n4339;
  assign n4341 = n889 & n4340;
  assign n4342 = n4338 & n4341;
  assign n4343 = n1931 & n4342;
  assign n4344 = n104 & n3481;
  assign n4345 = n701 & n4344;
  assign n4346 = n4343 & n4345;
  assign n4347 = n1281 & n4346;
  assign n4329 = n4144 ^ n4108;
  assign n4330 = ~n4141 & n4329;
  assign n4331 = n4330 ^ n4144;
  assign n4323 = n4139 ^ n4135;
  assign n4324 = ~n4136 & n4323;
  assign n4325 = n4324 ^ n4122;
  assign n4317 = n4134 ^ n2346;
  assign n4318 = n4126 & ~n4317;
  assign n4319 = n4318 ^ n2346;
  assign n4320 = n4319 ^ n2345;
  assign n4321 = ~n565 & ~n4320;
  assign n4310 = n573 & n2637;
  assign n4311 = n4310 ^ n2342;
  assign n4312 = n596 & n4311;
  assign n4313 = ~n2343 & ~n2488;
  assign n4314 = n2344 & n2492;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = ~n4312 & n4315;
  assign n4322 = n4321 ^ n4316;
  assign n4326 = n4325 ^ n4322;
  assign n4292 = n1108 & n3703;
  assign n4293 = ~n2320 & n2449;
  assign n4294 = ~n2360 & n2459;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = ~n4292 & n4295;
  assign n4297 = ~n595 & ~n4296;
  assign n4298 = n1108 & ~n3710;
  assign n4299 = n595 & n4295;
  assign n4300 = ~n4298 & n4299;
  assign n4301 = n2544 ^ n2317;
  assign n4302 = n4301 ^ n2544;
  assign n4303 = n618 & n1108;
  assign n4304 = n4303 ^ n2544;
  assign n4305 = ~n4302 & n4304;
  assign n4306 = n4305 ^ n2544;
  assign n4307 = n2382 & n4306;
  assign n4308 = ~n4300 & ~n4307;
  assign n4309 = ~n4297 & n4308;
  assign n4327 = n4326 ^ n4309;
  assign n4269 = ~n817 & n3163;
  assign n4270 = n4269 ^ n812;
  assign n4271 = n4270 ^ n3097;
  assign n4272 = n1451 & n4271;
  assign n4273 = ~n812 & n2425;
  assign n4274 = n3150 & n4273;
  assign n4275 = n4101 ^ n1100;
  assign n4276 = n4275 ^ n4101;
  assign n4277 = n3150 ^ n812;
  assign n4278 = n4277 ^ n4101;
  assign n4279 = n4276 & ~n4278;
  assign n4280 = n4279 ^ n4101;
  assign n4281 = ~n1451 & ~n4280;
  assign n4282 = n4281 ^ n816;
  assign n4283 = n4282 ^ n4281;
  assign n4284 = ~n3150 & n4096;
  assign n4285 = n2407 & n4094;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = n4286 ^ n4281;
  assign n4288 = ~n4283 & ~n4287;
  assign n4289 = n4288 ^ n4281;
  assign n4290 = ~n4274 & ~n4289;
  assign n4291 = ~n4272 & n4290;
  assign n4328 = n4327 ^ n4291;
  assign n4332 = n4331 ^ n4328;
  assign n4234 = n32 & n3676;
  assign n4235 = n3691 & ~n4234;
  assign n4236 = n2334 & n3643;
  assign n4237 = n2337 & ~n3116;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = n3853 ^ n3116;
  assign n4240 = n3643 ^ n3116;
  assign n4241 = n4239 & ~n4240;
  assign n4242 = n4241 ^ n3116;
  assign n4243 = n2815 ^ n2328;
  assign n4244 = ~n4242 & n4243;
  assign n4245 = n4238 & ~n4244;
  assign n4246 = n4245 ^ n2385;
  assign n4247 = n4246 ^ n4245;
  assign n4248 = n4245 ^ n3676;
  assign n4249 = n4248 ^ n4245;
  assign n4250 = n4247 & n4249;
  assign n4251 = n4250 ^ n4245;
  assign n4252 = n30 & n4251;
  assign n4253 = n4252 ^ n4245;
  assign n4254 = n4235 & n4253;
  assign n4255 = n2938 & ~n3691;
  assign n4256 = n3676 & n4255;
  assign n4257 = n30 & ~n4245;
  assign n4258 = ~n4256 & ~n4257;
  assign n4259 = ~n4254 & n4258;
  assign n4260 = n2385 ^ n30;
  assign n4261 = ~n3676 & ~n3691;
  assign n4262 = n4261 ^ n4245;
  assign n4263 = n4261 ^ n2385;
  assign n4264 = n4263 ^ n4261;
  assign n4265 = n4262 & ~n4264;
  assign n4266 = n4265 ^ n4261;
  assign n4267 = ~n4260 & n4266;
  assign n4268 = n4259 & ~n4267;
  assign n4333 = n4332 ^ n4268;
  assign n4206 = n3833 ^ x2;
  assign n4207 = n4206 ^ x2;
  assign n4208 = n3118 ^ x2;
  assign n4209 = ~n4207 & n4208;
  assign n4210 = n4209 ^ x2;
  assign n4211 = ~n3814 & n4210;
  assign n4212 = n4211 ^ x2;
  assign n4213 = n3180 & n4212;
  assign n4214 = ~x2 & ~x22;
  assign n4215 = n3188 & n4214;
  assign n4216 = x2 & x22;
  assign n4217 = n4216 ^ n3833;
  assign n4218 = n4216 ^ n3249;
  assign n4219 = n4218 ^ n3249;
  assign n4220 = n3249 ^ x1;
  assign n4221 = n4219 & ~n4220;
  assign n4222 = n4221 ^ n3249;
  assign n4223 = n4217 & ~n4222;
  assign n4224 = n4223 ^ n3833;
  assign n4225 = ~n4215 & ~n4224;
  assign n4226 = ~n4213 & n4225;
  assign n4227 = ~n3814 & ~n3833;
  assign n4228 = n4227 ^ x2;
  assign n4229 = n4228 ^ x2;
  assign n4230 = n3118 & n4229;
  assign n4231 = n4230 ^ x2;
  assign n4232 = n2325 & ~n4231;
  assign n4233 = n4226 & ~n4232;
  assign n4334 = n4333 ^ n4233;
  assign n4188 = ~n4145 & n4148;
  assign n4189 = n4153 ^ n4080;
  assign n4190 = ~n4081 & ~n4189;
  assign n4191 = n4190 ^ n4153;
  assign n4192 = n4188 & n4191;
  assign n4193 = n4061 & n4080;
  assign n4194 = ~n4188 & n4193;
  assign n4195 = ~n4153 & n4194;
  assign n4197 = ~n4061 & ~n4080;
  assign n4198 = n4153 & n4197;
  assign n4196 = n4145 & ~n4148;
  assign n4199 = n4198 ^ n4196;
  assign n4200 = n4199 ^ n4198;
  assign n4201 = n4198 ^ n4191;
  assign n4202 = n4200 & ~n4201;
  assign n4203 = n4202 ^ n4198;
  assign n4204 = ~n4195 & ~n4203;
  assign n4205 = ~n4192 & n4204;
  assign n4335 = n4334 ^ n4205;
  assign n4348 = n4347 ^ n4335;
  assign n4165 = ~n4021 & ~n4154;
  assign n4166 = ~n4004 & n4165;
  assign n4167 = ~n3797 & ~n3995;
  assign n4168 = n4166 & ~n4167;
  assign n4171 = n4154 ^ n4004;
  assign n4172 = n4154 ^ n4021;
  assign n4173 = n4171 & ~n4172;
  assign n4174 = n4173 ^ n4004;
  assign n4169 = n4021 & n4154;
  assign n4170 = n4004 & n4169;
  assign n4175 = n4174 ^ n4170;
  assign n4176 = n4175 ^ n4170;
  assign n4177 = n4170 ^ n3797;
  assign n4178 = n4177 ^ n4170;
  assign n4179 = ~n4176 & n4178;
  assign n4180 = n4179 ^ n4170;
  assign n4181 = ~n3987 & n4180;
  assign n4182 = n4181 ^ n4170;
  assign n4183 = ~n4168 & ~n4182;
  assign n4184 = ~n3797 & n4174;
  assign n4185 = n3995 & ~n4170;
  assign n4186 = n4184 & ~n4185;
  assign n4187 = n4183 & ~n4186;
  assign n4349 = n4348 ^ n4187;
  assign n4359 = n4348 ^ n4166;
  assign n4360 = n4359 ^ n4166;
  assign n4361 = n4172 ^ n4004;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = n4362 ^ n4166;
  assign n4364 = n3995 & n4363;
  assign n4350 = ~n4335 & n4347;
  assign n4351 = ~n4174 & ~n4350;
  assign n4352 = n4335 & ~n4347;
  assign n4353 = n3987 & ~n4166;
  assign n4354 = ~n4352 & n4353;
  assign n4355 = n4351 & n4354;
  assign n4356 = n3987 & n4170;
  assign n4357 = n4348 & n4356;
  assign n4358 = ~n4355 & ~n4357;
  assign n4365 = n4364 ^ n4358;
  assign n4469 = ~n4351 & ~n4352;
  assign n4470 = n4469 ^ n4364;
  assign n4464 = n4268 ^ n4233;
  assign n4465 = n4333 & ~n4464;
  assign n4466 = n4465 ^ n4233;
  assign n4459 = n4331 ^ n4327;
  assign n4460 = n4328 & n4459;
  assign n4461 = n4460 ^ n4291;
  assign n4454 = n4325 ^ n4309;
  assign n4455 = n4326 & ~n4454;
  assign n4456 = n4455 ^ n4309;
  assign n4446 = ~n565 & ~n4319;
  assign n4447 = n4446 ^ n2345;
  assign n4448 = n4446 ^ n4316;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = n4449 ^ n2345;
  assign n4451 = n4450 ^ n2344;
  assign n4452 = ~n565 & ~n4451;
  assign n4430 = n596 & n2422;
  assign n4431 = n2342 & ~n2488;
  assign n4432 = ~n2343 & n2492;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~n4430 & n4433;
  assign n4435 = ~n565 & ~n4434;
  assign n4436 = n596 & ~n2436;
  assign n4437 = n565 & n4433;
  assign n4438 = ~n4436 & n4437;
  assign n4439 = n2360 ^ n572;
  assign n4440 = n596 & n2421;
  assign n4441 = ~n4439 & n4440;
  assign n4442 = ~n4438 & ~n4441;
  assign n4443 = ~n4435 & n4442;
  assign n4444 = n4443 ^ n2327;
  assign n4416 = n2407 ^ n618;
  assign n4417 = n1108 & n4416;
  assign n4418 = n2384 & n4417;
  assign n4419 = n2317 & n2449;
  assign n4420 = ~n2320 & n2459;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = n595 & ~n4421;
  assign n4423 = ~n4418 & ~n4422;
  assign n4424 = n2413 & n2464;
  assign n4425 = n4423 & ~n4424;
  assign n4426 = n1108 & ~n2417;
  assign n4427 = ~n595 & n4421;
  assign n4428 = ~n4426 & n4427;
  assign n4429 = n4425 & ~n4428;
  assign n4445 = n4444 ^ n4429;
  assign n4453 = n4452 ^ n4445;
  assign n4457 = n4456 ^ n4453;
  assign n4402 = n1451 & n3845;
  assign n4403 = n2428 & ~n3097;
  assign n4404 = n2431 & ~n3150;
  assign n4405 = ~n4403 & ~n4404;
  assign n4406 = ~n4402 & n4405;
  assign n4407 = n812 & ~n4406;
  assign n4408 = n1451 & ~n3856;
  assign n4409 = ~n812 & n4405;
  assign n4410 = ~n4408 & n4409;
  assign n4411 = n1451 & n3144;
  assign n4412 = n3116 ^ n816;
  assign n4413 = n4411 & ~n4412;
  assign n4414 = ~n4410 & ~n4413;
  assign n4415 = ~n4407 & n4414;
  assign n4458 = n4457 ^ n4415;
  assign n4462 = n4461 ^ n4458;
  assign n4381 = ~n3815 & n3833;
  assign n4382 = n2385 & ~n4381;
  assign n4383 = n32 & ~n3643;
  assign n4384 = n2334 & ~n3691;
  assign n4385 = ~n2337 & ~n4384;
  assign n4386 = ~n4383 & ~n4385;
  assign n4387 = n2802 & ~n3691;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = n2329 & n3643;
  assign n4390 = n30 & ~n4389;
  assign n4391 = n4388 & n4390;
  assign n4392 = ~n4382 & n4391;
  assign n4393 = ~n3815 & ~n3833;
  assign n4394 = n2845 & n4393;
  assign n4395 = n3833 ^ n32;
  assign n4396 = n2385 & ~n4395;
  assign n4397 = n3815 & n4396;
  assign n4398 = ~n30 & ~n4388;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4394 & n4399;
  assign n4401 = ~n4392 & n4400;
  assign n4463 = n4462 ^ n4401;
  assign n4467 = n4466 ^ n4463;
  assign n4375 = ~n4198 & ~n4334;
  assign n4376 = ~n4195 & ~n4196;
  assign n4377 = ~n4375 & n4376;
  assign n4378 = ~n4188 & ~n4334;
  assign n4379 = n4191 & ~n4378;
  assign n4380 = ~n4377 & ~n4379;
  assign n4468 = n4467 ^ n4380;
  assign n4471 = n4470 ^ n4468;
  assign n4366 = n206 & n883;
  assign n4367 = n261 & ~n319;
  assign n4368 = n4366 & n4367;
  assign n4369 = n95 & ~n2389;
  assign n4370 = n406 & ~n4369;
  assign n4371 = n4368 & n4370;
  assign n4372 = n930 & n4371;
  assign n4373 = n2190 & n4372;
  assign n4374 = n735 & n4373;
  assign n4472 = n4471 ^ n4374;
  assign n4473 = n4472 ^ n4358;
  assign n4474 = n4473 ^ n4472;
  assign n4475 = n4472 ^ n3797;
  assign n4476 = n4474 & ~n4475;
  assign n4477 = n4476 ^ n4472;
  assign n4478 = n4365 & ~n4477;
  assign n4479 = n4478 ^ n4472;
  assign n4638 = ~n3797 & ~n4364;
  assign n4639 = ~n4374 & n4468;
  assign n4645 = ~n4469 & n4639;
  assign n4643 = n3797 & n4358;
  assign n4640 = n4374 & ~n4468;
  assign n4641 = ~n4469 & ~n4640;
  assign n4642 = ~n4639 & ~n4641;
  assign n4644 = n4643 ^ n4642;
  assign n4646 = n4645 ^ n4644;
  assign n4647 = n4646 ^ n4645;
  assign n4648 = n4468 ^ n4374;
  assign n4649 = n4648 ^ n4469;
  assign n4650 = n4649 ^ n4645;
  assign n4651 = n4650 ^ n4645;
  assign n4652 = n4647 & n4651;
  assign n4653 = n4652 ^ n4645;
  assign n4654 = ~n4638 & n4653;
  assign n4655 = n4654 ^ n4644;
  assign n4621 = ~n56 & n141;
  assign n4622 = n159 & ~n172;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = ~n403 & ~n4623;
  assign n4625 = ~n109 & n123;
  assign n4626 = ~n622 & n4625;
  assign n4627 = ~n297 & ~n4626;
  assign n4628 = n4624 & ~n4627;
  assign n4629 = n2052 & n4628;
  assign n4630 = n234 & ~n507;
  assign n4631 = n175 & n3524;
  assign n4632 = n4630 & n4631;
  assign n4633 = n4629 & n4632;
  assign n4634 = n3830 & n4633;
  assign n4635 = n3967 & n4634;
  assign n4636 = n3093 & n4635;
  assign n4615 = n4453 ^ n4415;
  assign n4616 = n4457 & n4615;
  assign n4617 = n4616 ^ n4415;
  assign n4581 = n2360 ^ n565;
  assign n4582 = n4581 ^ n2360;
  assign n4583 = n2826 & n4582;
  assign n4584 = n4583 ^ n2360;
  assign n4585 = ~n572 & ~n4584;
  assign n4586 = n4585 ^ n2360;
  assign n4587 = n2478 & ~n4586;
  assign n4588 = ~n572 & n2360;
  assign n4589 = n2342 & n2475;
  assign n4590 = ~n2487 & ~n4589;
  assign n4591 = ~n4588 & ~n4590;
  assign n4592 = ~n4587 & ~n4591;
  assign n4593 = n4592 ^ n565;
  assign n4594 = n596 & ~n2842;
  assign n4595 = n4594 ^ n565;
  assign n4596 = n565 & n596;
  assign n4597 = n2846 & n4596;
  assign n4598 = n2320 ^ n572;
  assign n4599 = n596 & n2841;
  assign n4600 = n4598 & n4599;
  assign n4601 = ~n4597 & ~n4600;
  assign n4602 = n4601 ^ n565;
  assign n4603 = ~n565 & ~n4602;
  assign n4604 = n4603 ^ n565;
  assign n4605 = ~n4595 & ~n4604;
  assign n4606 = n4605 ^ n4603;
  assign n4607 = n4606 ^ n565;
  assign n4608 = n4607 ^ n4601;
  assign n4609 = n4593 & ~n4608;
  assign n4610 = n4609 ^ n4601;
  assign n4567 = ~n2327 & n4443;
  assign n4568 = n2344 & n4567;
  assign n4569 = ~n565 & ~n2343;
  assign n4570 = ~n4568 & n4569;
  assign n4571 = n2327 & ~n4443;
  assign n4572 = ~n2344 & n4571;
  assign n4573 = n4570 & ~n4572;
  assign n4574 = n565 & n4571;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = n2343 & n4572;
  assign n4534 = ~n565 & n2344;
  assign n4577 = n2343 & n4534;
  assign n4578 = n4567 & n4577;
  assign n4579 = ~n4576 & ~n4578;
  assign n4580 = n4575 & n4579;
  assign n4611 = n4610 ^ n4580;
  assign n4545 = ~n2407 & n2449;
  assign n4546 = n2317 & n2459;
  assign n4547 = ~n4545 & ~n4546;
  assign n4548 = n595 & n4547;
  assign n4549 = n3150 ^ n618;
  assign n4550 = n4549 ^ n3150;
  assign n4551 = n3185 ^ n3150;
  assign n4552 = ~n4550 & n4551;
  assign n4553 = n4552 ^ n3150;
  assign n4554 = n1108 & ~n4553;
  assign n4555 = n4548 & ~n4554;
  assign n4556 = n618 & n3184;
  assign n4557 = ~n595 & ~n3150;
  assign n4558 = n1108 & n4557;
  assign n4559 = ~n4556 & n4558;
  assign n4560 = ~n595 & ~n4547;
  assign n4561 = ~n595 & n4303;
  assign n4562 = n3150 & n4561;
  assign n4563 = n3184 & n4562;
  assign n4564 = ~n4560 & ~n4563;
  assign n4565 = ~n4559 & n4564;
  assign n4566 = ~n4555 & n4565;
  assign n4612 = n4611 ^ n4566;
  assign n4535 = n4429 & n4444;
  assign n4536 = ~n4534 & n4535;
  assign n4537 = n4444 ^ n2344;
  assign n4538 = ~n4450 & n4537;
  assign n4539 = ~n4429 & ~n4538;
  assign n4540 = n2344 & ~n4444;
  assign n4541 = n4450 & ~n4540;
  assign n4542 = ~n565 & ~n4541;
  assign n4543 = ~n4539 & n4542;
  assign n4544 = ~n4536 & ~n4543;
  assign n4613 = n4612 ^ n4544;
  assign n4519 = n3643 & ~n3655;
  assign n4520 = n1451 & n4519;
  assign n4521 = n2428 & ~n3116;
  assign n4522 = n2431 & ~n3097;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = ~n4520 & n4523;
  assign n4525 = ~n812 & ~n4524;
  assign n4526 = n1451 & ~n4047;
  assign n4527 = n812 & n4523;
  assign n4528 = ~n4526 & n4527;
  assign n4529 = n3643 ^ n816;
  assign n4530 = n1451 & ~n4529;
  assign n4531 = n3655 & n4530;
  assign n4532 = ~n4528 & ~n4531;
  assign n4533 = ~n4525 & n4532;
  assign n4614 = n4613 ^ n4533;
  assign n4618 = n4617 ^ n4614;
  assign n4502 = ~n2803 & ~n3833;
  assign n4503 = n2337 & ~n3691;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = ~n30 & ~n4504;
  assign n4506 = n30 & ~n4502;
  assign n4507 = ~n32 & ~n2327;
  assign n4508 = ~n3691 & n4507;
  assign n4509 = n4506 & ~n4508;
  assign n4510 = ~n2385 & ~n4509;
  assign n4511 = ~n32 & n2385;
  assign n4512 = n4511 ^ n4506;
  assign n4513 = n4511 ^ n4066;
  assign n4514 = n4513 ^ n4511;
  assign n4515 = ~n4512 & ~n4514;
  assign n4516 = n4515 ^ n4511;
  assign n4517 = ~n4510 & ~n4516;
  assign n4518 = ~n4505 & ~n4517;
  assign n4619 = n4618 ^ n4518;
  assign n4480 = ~n4401 & ~n4466;
  assign n4481 = n4380 & ~n4480;
  assign n4482 = n4458 & ~n4461;
  assign n4483 = ~n4458 & n4461;
  assign n4484 = n4401 & ~n4483;
  assign n4485 = n4466 & n4484;
  assign n4486 = ~n4482 & ~n4485;
  assign n4487 = n4481 & ~n4486;
  assign n4489 = n4458 ^ n4401;
  assign n4490 = n4489 ^ n4461;
  assign n4491 = n4482 & ~n4490;
  assign n4492 = n4491 ^ n4490;
  assign n4493 = ~n4466 & ~n4492;
  assign n4488 = ~n4401 & n4483;
  assign n4494 = n4493 ^ n4488;
  assign n4495 = ~n4380 & n4494;
  assign n4496 = n4401 & n4482;
  assign n4497 = n4496 ^ n4488;
  assign n4498 = n4466 & n4497;
  assign n4499 = n4498 ^ n4488;
  assign n4500 = ~n4495 & ~n4499;
  assign n4501 = ~n4487 & n4500;
  assign n4620 = n4619 ^ n4501;
  assign n4637 = n4636 ^ n4620;
  assign n4656 = n4655 ^ n4637;
  assign n4793 = n4642 ^ n4620;
  assign n4794 = n4637 & ~n4793;
  assign n4795 = n4794 ^ n4642;
  assign n4774 = ~n45 & ~n167;
  assign n4775 = n101 & ~n4774;
  assign n4776 = ~n823 & ~n4775;
  assign n4777 = n3959 & ~n4776;
  assign n4778 = n3818 & n4777;
  assign n4779 = n175 & ~n197;
  assign n4780 = n1923 & n4779;
  assign n4781 = n2251 & n4780;
  assign n4782 = n4778 & n4781;
  assign n4783 = ~n111 & ~n525;
  assign n4784 = n2077 & n4783;
  assign n4785 = n688 & n4784;
  assign n4786 = ~n105 & ~n472;
  assign n4787 = n3106 & n4786;
  assign n4788 = n4785 & n4787;
  assign n4789 = n4782 & n4788;
  assign n4790 = n2180 & n4789;
  assign n4791 = n3522 & n4790;
  assign n4768 = n4544 ^ n4533;
  assign n4769 = ~n4613 & n4768;
  assign n4770 = n4769 ^ n4533;
  assign n4763 = n4580 ^ n4566;
  assign n4764 = ~n4611 & n4763;
  assign n4765 = n4764 ^ n4566;
  assign n4744 = ~n565 & ~n2320;
  assign n4745 = n2487 & n4744;
  assign n4746 = n2490 & n4588;
  assign n4747 = ~n565 & n2360;
  assign n4748 = n2301 & ~n4747;
  assign n4749 = ~n4746 & ~n4748;
  assign n4750 = ~n4745 & n4749;
  assign n4751 = n2320 ^ n565;
  assign n4752 = n565 & n611;
  assign n4753 = ~n2479 & ~n4752;
  assign n4754 = ~n4751 & ~n4753;
  assign n4755 = n4750 & ~n4754;
  assign n4756 = n573 & ~n2382;
  assign n4757 = n4756 ^ n572;
  assign n4758 = n4757 ^ n2317;
  assign n4759 = n596 & n4758;
  assign n4760 = n4755 & ~n4759;
  assign n4731 = n4568 & n4569;
  assign n4732 = ~n4576 & ~n4731;
  assign n4733 = ~n2342 & ~n4732;
  assign n4734 = ~n2343 & n2344;
  assign n4735 = n4443 & n4734;
  assign n4736 = ~n565 & n2342;
  assign n4737 = ~n4735 & n4736;
  assign n4738 = ~n4576 & n4737;
  assign n4739 = n2327 & n4569;
  assign n4740 = n2342 & n4739;
  assign n4741 = ~n4574 & ~n4740;
  assign n4742 = ~n4738 & n4741;
  assign n4743 = ~n4733 & n4742;
  assign n4761 = n4760 ^ n4743;
  assign n4716 = n1108 & ~n3097;
  assign n4717 = ~n3163 & n4716;
  assign n4718 = n2449 & ~n3150;
  assign n4719 = ~n2407 & n2459;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4717 & n4720;
  assign n4722 = ~n595 & ~n4721;
  assign n4723 = n1108 & n3163;
  assign n4726 = n3097 ^ n618;
  assign n4724 = n595 & n4720;
  assign n4725 = ~n4716 & n4724;
  assign n4727 = n4726 ^ n4725;
  assign n4728 = n4723 & ~n4727;
  assign n4729 = n4728 ^ n4725;
  assign n4730 = ~n4722 & ~n4729;
  assign n4762 = n4761 ^ n4730;
  assign n4766 = n4765 ^ n4762;
  assign n4701 = n1451 & n4261;
  assign n4702 = n2428 & n3643;
  assign n4703 = n2431 & ~n3116;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = ~n4701 & n4704;
  assign n4706 = ~n812 & ~n4705;
  assign n4707 = ~n3676 & n3691;
  assign n4708 = n1451 & ~n4707;
  assign n4709 = n812 & n4704;
  assign n4710 = ~n4708 & n4709;
  assign n4711 = n3691 ^ n816;
  assign n4712 = n1451 & n4711;
  assign n4713 = n3676 & n4712;
  assign n4714 = ~n4710 & ~n4713;
  assign n4715 = ~n4706 & n4714;
  assign n4767 = n4766 ^ n4715;
  assign n4771 = n4770 ^ n4767;
  assign n4697 = n4614 ^ n4518;
  assign n4698 = n4618 & n4697;
  assign n4699 = n4698 ^ n4518;
  assign n4684 = n3814 ^ n30;
  assign n4685 = n4684 ^ n30;
  assign n4686 = ~n32 & ~n3833;
  assign n4687 = n4686 ^ n30;
  assign n4688 = ~n4685 & ~n4687;
  assign n4689 = n4688 ^ n30;
  assign n4690 = ~n2333 & ~n4689;
  assign n4691 = n2328 ^ n32;
  assign n4692 = n2328 ^ n30;
  assign n4693 = n4691 & ~n4692;
  assign n4694 = ~n3833 & n4693;
  assign n4695 = n4694 ^ n30;
  assign n4696 = ~n4690 & n4695;
  assign n4700 = n4699 ^ n4696;
  assign n4772 = n4771 ^ n4700;
  assign n4672 = ~n4485 & n4619;
  assign n4673 = n4380 & ~n4672;
  assign n4674 = ~n4480 & ~n4619;
  assign n4675 = ~n4482 & ~n4674;
  assign n4676 = ~n4673 & n4675;
  assign n4677 = ~n4483 & ~n4619;
  assign n4678 = n4466 ^ n4380;
  assign n4679 = n4401 ^ n4380;
  assign n4680 = n4678 & n4679;
  assign n4681 = n4680 ^ n4380;
  assign n4682 = ~n4677 & ~n4681;
  assign n4683 = ~n4676 & ~n4682;
  assign n4773 = n4772 ^ n4683;
  assign n4792 = n4791 ^ n4773;
  assign n4796 = n4795 ^ n4792;
  assign n4658 = n4469 & n4640;
  assign n4657 = ~n4642 & ~n4645;
  assign n4659 = n4658 ^ n4657;
  assign n4660 = n4637 & n4659;
  assign n4661 = n4660 ^ n4657;
  assign n4662 = ~n4358 & n4661;
  assign n4663 = n3797 & ~n4662;
  assign n4664 = ~n4637 & n4641;
  assign n4665 = n4364 & ~n4658;
  assign n4666 = ~n4664 & n4665;
  assign n4667 = n4637 ^ n4469;
  assign n4668 = ~n4639 & n4667;
  assign n4669 = n4668 ^ n4469;
  assign n4670 = n4666 & ~n4669;
  assign n4671 = ~n4663 & ~n4670;
  assign n4797 = n4796 ^ n4671;
  assign n4913 = n4795 ^ n4773;
  assign n4914 = ~n4792 & n4913;
  assign n4915 = n4914 ^ n4795;
  assign n4893 = ~n4767 & n4770;
  assign n4894 = ~n4696 & n4893;
  assign n4895 = n4767 & ~n4770;
  assign n4896 = n4696 & n4895;
  assign n4897 = ~n4894 & ~n4896;
  assign n4898 = n4700 & ~n4897;
  assign n4899 = ~n4696 & ~n4895;
  assign n4900 = ~n4893 & ~n4899;
  assign n4901 = ~n4699 & ~n4894;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = n4902 ^ n4683;
  assign n4904 = n4903 ^ n4902;
  assign n4905 = ~n4699 & n4900;
  assign n4906 = ~n4896 & ~n4905;
  assign n4907 = n4906 ^ n4902;
  assign n4908 = ~n4904 & ~n4907;
  assign n4909 = n4908 ^ n4902;
  assign n4910 = ~n4898 & ~n4909;
  assign n4878 = n1451 & n4393;
  assign n4879 = n2431 & n3643;
  assign n4880 = n2428 & ~n3691;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~n4878 & n4881;
  assign n4883 = n812 & ~n4882;
  assign n4884 = n1451 & ~n4381;
  assign n4885 = ~n812 & n4881;
  assign n4886 = ~n4884 & n4885;
  assign n4887 = n3833 ^ n816;
  assign n4888 = n1451 & ~n4887;
  assign n4889 = n3815 & n4888;
  assign n4890 = ~n4886 & ~n4889;
  assign n4891 = ~n4883 & n4890;
  assign n4874 = n4762 ^ n4715;
  assign n4875 = n4766 & ~n4874;
  assign n4876 = n4875 ^ n4715;
  assign n4844 = ~n618 & n3144;
  assign n4845 = ~n3116 & ~n4844;
  assign n4846 = n2449 & ~n3097;
  assign n4847 = n2459 & ~n3150;
  assign n4848 = ~n4846 & ~n4847;
  assign n4849 = n4848 ^ n1108;
  assign n4850 = n4849 ^ n1108;
  assign n4851 = n3144 ^ n1108;
  assign n4852 = n4851 ^ n1108;
  assign n4853 = n4850 & n4852;
  assign n4854 = n4853 ^ n1108;
  assign n4855 = ~n595 & n4854;
  assign n4856 = n4855 ^ n1108;
  assign n4857 = n4845 & n4856;
  assign n4858 = n4848 ^ n595;
  assign n4859 = n1108 & ~n3856;
  assign n4860 = n4859 ^ n595;
  assign n4861 = n2544 & n3116;
  assign n4862 = n3144 & n4861;
  assign n4863 = n4862 ^ n595;
  assign n4864 = ~n595 & n4863;
  assign n4865 = n4864 ^ n595;
  assign n4866 = ~n4860 & ~n4865;
  assign n4867 = n4866 ^ n4864;
  assign n4868 = n4867 ^ n595;
  assign n4869 = n4868 ^ n4862;
  assign n4870 = n4858 & n4869;
  assign n4871 = n4870 ^ n4862;
  assign n4872 = ~n4857 & ~n4871;
  assign n4840 = n4743 ^ n4730;
  assign n4841 = n4761 & n4840;
  assign n4842 = n4841 ^ n4730;
  assign n4813 = n2317 & ~n2488;
  assign n4814 = ~n2320 & n2492;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = n573 & n2384;
  assign n4817 = n4816 ^ n2407;
  assign n4818 = n596 & ~n4817;
  assign n4819 = n4815 & ~n4818;
  assign n4820 = ~n2327 & n2342;
  assign n4821 = n4735 & n4820;
  assign n4822 = n2360 & n4821;
  assign n4823 = n565 & ~n4571;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = n4819 & ~n4824;
  assign n4826 = ~n4534 & ~n4569;
  assign n4827 = ~n4736 & n4826;
  assign n4828 = ~n4443 & n4827;
  assign n4829 = n2327 & n4828;
  assign n4830 = ~n2360 & ~n4829;
  assign n4831 = n4830 ^ n4819;
  assign n4832 = n4831 ^ n4830;
  assign n4833 = ~n4747 & ~n4829;
  assign n4834 = n4833 ^ n4830;
  assign n4835 = ~n4832 & ~n4834;
  assign n4836 = n4835 ^ n4830;
  assign n4837 = ~n4821 & n4836;
  assign n4838 = ~n4825 & ~n4837;
  assign n4839 = n4838 ^ n30;
  assign n4843 = n4842 ^ n4839;
  assign n4873 = n4872 ^ n4843;
  assign n4877 = n4876 ^ n4873;
  assign n4892 = n4891 ^ n4877;
  assign n4911 = n4910 ^ n4892;
  assign n4803 = ~n166 & ~n3470;
  assign n4804 = ~n270 & n451;
  assign n4805 = n683 & ~n4804;
  assign n4806 = ~n551 & ~n719;
  assign n4807 = n4805 & ~n4806;
  assign n4808 = n3052 & n4624;
  assign n4809 = n4807 & n4808;
  assign n4810 = n4782 & n4809;
  assign n4811 = ~n4803 & n4810;
  assign n4812 = n1993 & n4811;
  assign n4912 = n4911 ^ n4812;
  assign n4916 = n4915 ^ n4912;
  assign n4798 = n4662 & ~n4670;
  assign n4799 = n4796 & n4798;
  assign n4800 = n4670 & ~n4796;
  assign n4801 = ~n3797 & ~n4800;
  assign n4802 = ~n4799 & ~n4801;
  assign n4917 = n4916 ^ n4802;
  assign n5037 = n60 & ~n535;
  assign n5038 = n372 & ~n5037;
  assign n5039 = n71 & n2389;
  assign n5040 = n172 & ~n5039;
  assign n5041 = n5038 & ~n5040;
  assign n5042 = n1905 & n5041;
  assign n5043 = n3523 & n5042;
  assign n5044 = n138 & n2077;
  assign n5045 = n2233 & n3082;
  assign n5046 = n5044 & n5045;
  assign n5047 = n110 & ~n159;
  assign n5048 = n59 & ~n120;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = ~n2123 & n5049;
  assign n5051 = n921 & n5050;
  assign n5052 = n5046 & n5051;
  assign n5053 = n5043 & n5052;
  assign n5054 = n3462 & n5053;
  assign n5031 = n4872 ^ n4839;
  assign n5032 = ~n4843 & ~n5031;
  assign n5033 = n5032 ^ n4842;
  assign n5015 = n2428 & ~n3833;
  assign n5016 = n2431 & ~n3691;
  assign n5017 = ~n5015 & ~n5016;
  assign n5018 = n5017 ^ n812;
  assign n5019 = n5018 ^ n816;
  assign n5020 = n5018 ^ n5017;
  assign n5021 = n1451 & n4066;
  assign n5022 = n5021 ^ n5017;
  assign n5023 = ~n5017 & ~n5022;
  assign n5024 = n5023 ^ n5017;
  assign n5025 = ~n5020 & ~n5024;
  assign n5026 = n5025 ^ n5023;
  assign n5027 = n5026 ^ n5017;
  assign n5028 = n5027 ^ n5021;
  assign n5029 = n5019 & ~n5028;
  assign n5030 = n5029 ^ n5018;
  assign n5034 = n5033 ^ n5030;
  assign n5011 = n4891 ^ n4873;
  assign n5012 = n4877 & n5011;
  assign n5013 = n5012 ^ n4876;
  assign n4983 = n4735 & n4736;
  assign n4984 = n2327 & ~n4828;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = n565 & ~n4819;
  assign n4987 = ~n4985 & n4986;
  assign n4988 = ~n2327 & ~n2360;
  assign n4989 = n4819 & ~n4988;
  assign n4990 = ~n2360 & ~n4985;
  assign n4991 = ~n4989 & ~n4990;
  assign n4992 = ~n565 & ~n4991;
  assign n4993 = ~n4983 & ~n4986;
  assign n4994 = ~n2327 & ~n4993;
  assign n4995 = ~n4992 & ~n4994;
  assign n4996 = n4995 ^ n30;
  assign n4997 = n4996 ^ n4995;
  assign n4998 = n2360 & ~n4985;
  assign n4999 = ~n4986 & ~n4998;
  assign n5000 = n2327 & ~n4999;
  assign n5001 = ~n565 & n4988;
  assign n5002 = n4985 & ~n5001;
  assign n5003 = n4819 & ~n5002;
  assign n5004 = ~n5000 & ~n5003;
  assign n5005 = n5004 ^ n4995;
  assign n5006 = ~n4997 & n5005;
  assign n5007 = n5006 ^ n4995;
  assign n5008 = ~n4987 & n5007;
  assign n4972 = n2327 ^ n30;
  assign n4973 = n2327 ^ n565;
  assign n4974 = n4973 ^ n2327;
  assign n4975 = n2360 ^ n2327;
  assign n4976 = n4975 ^ n2327;
  assign n4977 = ~n4974 & ~n4976;
  assign n4978 = n4977 ^ n2327;
  assign n4979 = n4972 & n4978;
  assign n4980 = n4979 ^ n30;
  assign n4981 = n4980 ^ n4744;
  assign n4957 = n596 & ~n3150;
  assign n4958 = ~n3184 & n4957;
  assign n4959 = ~n2407 & ~n2488;
  assign n4960 = n2317 & n2492;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = ~n4958 & n4961;
  assign n4963 = ~n565 & ~n4962;
  assign n4964 = n3150 ^ n572;
  assign n4965 = n596 & ~n4964;
  assign n4966 = n3184 & n4965;
  assign n4967 = ~n4963 & ~n4966;
  assign n4968 = n596 & ~n3547;
  assign n4969 = n565 & n4961;
  assign n4970 = ~n4968 & n4969;
  assign n4971 = n4967 & ~n4970;
  assign n4982 = n4981 ^ n4971;
  assign n5009 = n5008 ^ n4982;
  assign n4938 = ~n618 & n3643;
  assign n4939 = ~n4519 & ~n4938;
  assign n4940 = n1108 & ~n4939;
  assign n4941 = n2449 & ~n3116;
  assign n4942 = n2459 & ~n3097;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~n4940 & n4943;
  assign n4945 = ~n595 & ~n4944;
  assign n4946 = n595 & n4943;
  assign n4947 = n3643 ^ n618;
  assign n4948 = n4947 ^ n3643;
  assign n4949 = n3656 ^ n3643;
  assign n4950 = ~n4948 & n4949;
  assign n4951 = n4950 ^ n3643;
  assign n4952 = n1108 & n4951;
  assign n4953 = n4946 & ~n4952;
  assign n4954 = n4050 & n4561;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = ~n4945 & n4955;
  assign n5010 = n5009 ^ n4956;
  assign n5014 = n5013 ^ n5010;
  assign n5035 = n5034 ^ n5014;
  assign n4925 = ~n4892 & ~n4895;
  assign n4926 = n4699 ^ n4683;
  assign n4927 = n4700 & n4926;
  assign n4928 = n4927 ^ n4683;
  assign n4929 = ~n4925 & ~n4928;
  assign n4930 = n4699 & n4899;
  assign n4931 = n4892 & ~n4930;
  assign n4932 = n4683 & ~n4931;
  assign n4933 = n4696 & ~n4699;
  assign n4934 = ~n4892 & ~n4933;
  assign n4935 = ~n4893 & ~n4934;
  assign n4936 = ~n4932 & n4935;
  assign n4937 = ~n4929 & ~n4936;
  assign n5036 = n5035 ^ n4937;
  assign n5055 = n5054 ^ n5036;
  assign n4922 = n4915 ^ n4911;
  assign n4923 = n4912 & ~n4922;
  assign n4924 = n4923 ^ n4915;
  assign n5056 = n5055 ^ n4924;
  assign n4918 = n4799 & ~n4916;
  assign n4919 = n3797 & ~n4918;
  assign n4920 = n4800 & n4916;
  assign n4921 = ~n4919 & ~n4920;
  assign n5057 = n5056 ^ n4921;
  assign n5152 = ~n3797 & ~n4920;
  assign n5153 = n5152 ^ n4919;
  assign n5154 = n5054 ^ n4919;
  assign n5155 = n5154 ^ n4919;
  assign n5156 = n5153 & n5155;
  assign n5157 = n5156 ^ n4919;
  assign n5158 = n5055 & n5157;
  assign n5159 = n5036 & ~n5152;
  assign n5160 = n5159 ^ n5054;
  assign n5161 = ~n5154 & ~n5160;
  assign n5162 = n5161 ^ n5054;
  assign n5163 = n5162 ^ n4924;
  assign n5164 = n5163 ^ n5162;
  assign n5165 = ~n5036 & n5054;
  assign n5166 = ~n4919 & n5165;
  assign n5167 = n5036 & ~n5054;
  assign n5168 = n5152 & ~n5167;
  assign n5169 = ~n5166 & ~n5168;
  assign n5170 = n5169 ^ n5162;
  assign n5171 = n5164 & n5170;
  assign n5172 = n5171 ^ n5162;
  assign n5173 = ~n5158 & n5172;
  assign n5142 = ~n426 & n2036;
  assign n5143 = ~n126 & ~n659;
  assign n5144 = n642 & n5143;
  assign n5145 = n5142 & n5144;
  assign n5146 = n3955 & n5145;
  assign n5147 = n685 & n4787;
  assign n5148 = n5146 & n5147;
  assign n5149 = n3529 & n5148;
  assign n5150 = n2254 & n5149;
  assign n5119 = n3814 ^ n812;
  assign n5120 = n5119 ^ n812;
  assign n5121 = n816 & ~n3833;
  assign n5122 = n5121 ^ n812;
  assign n5123 = ~n5120 & ~n5122;
  assign n5124 = n5123 ^ n812;
  assign n5125 = ~n2424 & ~n5124;
  assign n5126 = ~n812 & n816;
  assign n5127 = ~n2425 & ~n5126;
  assign n5128 = n5127 ^ n812;
  assign n5129 = n3833 ^ n812;
  assign n5130 = n5129 ^ n812;
  assign n5131 = n5128 & ~n5130;
  assign n5132 = n5131 ^ n812;
  assign n5133 = n5125 ^ n2746;
  assign n5134 = n5132 & ~n5133;
  assign n5135 = n5134 ^ n2746;
  assign n5136 = ~n5125 & n5135;
  assign n5137 = n5136 ^ n5125;
  assign n5138 = n5137 ^ n5125;
  assign n5116 = n5008 ^ n4956;
  assign n5117 = n5009 & n5116;
  assign n5118 = n5117 ^ n4956;
  assign n5139 = n5138 ^ n5118;
  assign n5113 = ~n565 & n2383;
  assign n5094 = ~n2407 & n2504;
  assign n5095 = n611 & ~n5094;
  assign n5096 = n2479 & ~n3150;
  assign n5097 = n5096 ^ n2478;
  assign n5098 = ~n5095 & ~n5097;
  assign n5099 = n3150 ^ n2407;
  assign n5100 = n5099 ^ n3150;
  assign n5101 = n3150 ^ n565;
  assign n5102 = n5101 ^ n3150;
  assign n5103 = ~n5100 & n5102;
  assign n5104 = n5103 ^ n3150;
  assign n5105 = n595 & ~n5104;
  assign n5106 = n5105 ^ n3150;
  assign n5107 = ~n572 & ~n5106;
  assign n5108 = ~n5098 & ~n5107;
  assign n5109 = n573 & n3163;
  assign n5110 = n5109 ^ n3097;
  assign n5111 = n596 & n5110;
  assign n5112 = ~n5108 & ~n5111;
  assign n5114 = n5113 ^ n5112;
  assign n5089 = n4971 ^ n4744;
  assign n5090 = n4980 ^ n4971;
  assign n5091 = ~n5089 & n5090;
  assign n5092 = n5091 ^ n4744;
  assign n5075 = n1108 & n4261;
  assign n5076 = n2449 & n3643;
  assign n5077 = n2459 & ~n3116;
  assign n5078 = ~n5076 & ~n5077;
  assign n5079 = ~n5075 & n5078;
  assign n5080 = ~n595 & ~n5079;
  assign n5081 = n1108 & ~n4707;
  assign n5082 = n595 & n5078;
  assign n5083 = ~n5081 & n5082;
  assign n5084 = n3691 ^ n618;
  assign n5085 = n1108 & ~n5084;
  assign n5086 = n3676 & n5085;
  assign n5087 = ~n5083 & ~n5086;
  assign n5088 = ~n5080 & n5087;
  assign n5093 = n5092 ^ n5088;
  assign n5115 = n5114 ^ n5093;
  assign n5140 = n5139 ^ n5115;
  assign n5058 = ~n5010 & n5013;
  assign n5059 = ~n5030 & ~n5033;
  assign n5065 = ~n5058 & n5059;
  assign n5061 = n5010 & ~n5013;
  assign n5062 = n5030 & n5033;
  assign n5066 = n5061 & ~n5062;
  assign n5067 = ~n5065 & ~n5066;
  assign n5060 = n5058 & ~n5059;
  assign n5063 = ~n5061 & n5062;
  assign n5064 = ~n5060 & ~n5063;
  assign n5068 = n5067 ^ n5064;
  assign n5069 = ~n4937 & n5068;
  assign n5070 = n5069 ^ n5064;
  assign n5071 = n5030 ^ n5010;
  assign n5072 = ~n5034 & n5071;
  assign n5073 = n5014 & n5072;
  assign n5074 = n5070 & ~n5073;
  assign n5141 = n5140 ^ n5074;
  assign n5151 = n5150 ^ n5141;
  assign n5174 = n5173 ^ n5151;
  assign n5272 = n5167 ^ n5150;
  assign n5273 = n5272 ^ n5150;
  assign n5179 = ~n4924 & ~n5165;
  assign n5274 = n5179 ^ n5150;
  assign n5275 = n5274 ^ n5150;
  assign n5276 = ~n5273 & ~n5275;
  assign n5277 = n5276 ^ n5150;
  assign n5278 = ~n5151 & ~n5277;
  assign n5279 = n5278 ^ n5141;
  assign n5263 = n86 & ~n408;
  assign n5264 = n3454 & ~n5263;
  assign n5265 = ~n549 & ~n2198;
  assign n5266 = n5264 & n5265;
  assign n5267 = n3964 & n5266;
  assign n5268 = n448 & n5267;
  assign n5269 = n1032 & n3482;
  assign n5270 = n5268 & n5269;
  assign n5257 = n5114 ^ n5092;
  assign n5258 = n5093 & ~n5257;
  assign n5259 = n5258 ^ n5088;
  assign n5234 = n573 & ~n3144;
  assign n5235 = n5234 ^ n572;
  assign n5236 = n5235 ^ n3116;
  assign n5237 = n596 & n5236;
  assign n5238 = ~n565 & n2478;
  assign n5239 = n3097 & n5238;
  assign n5240 = n3097 ^ n565;
  assign n5241 = n611 & n5240;
  assign n5242 = n2490 & n3150;
  assign n5243 = n5242 ^ n2478;
  assign n5244 = ~n5241 & ~n5243;
  assign n5245 = n5244 ^ n572;
  assign n5246 = n5245 ^ n5244;
  assign n5247 = n2490 & ~n3097;
  assign n5248 = ~n565 & n3150;
  assign n5249 = n611 & n5248;
  assign n5250 = ~n5247 & ~n5249;
  assign n5251 = n5250 ^ n5244;
  assign n5252 = n5246 & n5251;
  assign n5253 = n5252 ^ n5244;
  assign n5254 = ~n5239 & n5253;
  assign n5255 = ~n5237 & n5254;
  assign n5227 = n5112 ^ n565;
  assign n5228 = n5227 ^ n2317;
  assign n5229 = n5112 ^ n2320;
  assign n5230 = ~n2383 & ~n5229;
  assign n5231 = ~n5228 & n5230;
  assign n5232 = n5231 ^ n5227;
  assign n5224 = n2407 ^ n2320;
  assign n5225 = ~n565 & n5224;
  assign n5226 = n5225 ^ n812;
  assign n5233 = n5232 ^ n5226;
  assign n5256 = n5255 ^ n5233;
  assign n5260 = n5259 ^ n5256;
  assign n5220 = n5118 ^ n5115;
  assign n5221 = n5139 & n5220;
  assign n5222 = n5221 ^ n5115;
  assign n5206 = n1108 & ~n4381;
  assign n5207 = n2459 & n3643;
  assign n5208 = n2449 & ~n3691;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = ~n595 & n5209;
  assign n5211 = ~n5206 & n5210;
  assign n5212 = n2464 & n4393;
  assign n5213 = n3833 ^ n618;
  assign n5214 = n1108 & n5213;
  assign n5215 = n3815 & n5214;
  assign n5216 = n595 & ~n5209;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5212 & n5217;
  assign n5219 = ~n5211 & n5218;
  assign n5223 = n5222 ^ n5219;
  assign n5261 = n5260 ^ n5223;
  assign n5196 = ~n5059 & ~n5140;
  assign n5197 = ~n5060 & ~n5196;
  assign n5198 = ~n5061 & ~n5140;
  assign n5199 = ~n5063 & ~n5198;
  assign n5200 = n5197 & n5199;
  assign n5201 = n4937 & ~n5200;
  assign n5202 = n5062 & ~n5197;
  assign n5203 = ~n5065 & n5198;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n5201 & n5204;
  assign n5262 = n5261 ^ n5205;
  assign n5271 = n5270 ^ n5262;
  assign n5280 = n5279 ^ n5271;
  assign n5175 = n4924 & n5055;
  assign n5176 = n4920 & ~n5175;
  assign n5177 = n5167 ^ n5151;
  assign n5178 = n5177 ^ n5167;
  assign n5180 = n5179 ^ n5167;
  assign n5181 = ~n5178 & ~n5180;
  assign n5182 = n5181 ^ n5167;
  assign n5183 = n5176 & n5182;
  assign n5184 = ~n3797 & ~n5183;
  assign n5185 = n5151 & ~n5165;
  assign n5186 = n4918 & ~n5185;
  assign n5187 = n5165 ^ n4924;
  assign n5188 = n5187 ^ n5165;
  assign n5189 = n5165 ^ n5151;
  assign n5190 = n5188 & n5189;
  assign n5191 = n5190 ^ n5165;
  assign n5192 = ~n5167 & ~n5191;
  assign n5193 = n5192 ^ n4924;
  assign n5194 = n5186 & n5193;
  assign n5195 = ~n5184 & ~n5194;
  assign n5281 = n5280 ^ n5195;
  assign n5359 = n5279 ^ n5262;
  assign n5360 = ~n5271 & ~n5359;
  assign n5361 = n5360 ^ n5279;
  assign n5338 = ~n5256 & ~n5259;
  assign n5339 = n5219 & n5338;
  assign n5340 = n5256 & n5259;
  assign n5341 = ~n5219 & n5340;
  assign n5342 = ~n5339 & ~n5341;
  assign n5343 = n5223 & ~n5342;
  assign n5344 = n5259 ^ n5219;
  assign n5345 = ~n5260 & ~n5344;
  assign n5346 = n5345 ^ n5219;
  assign n5347 = ~n5222 & n5346;
  assign n5348 = ~n5339 & ~n5347;
  assign n5349 = n5348 ^ n5205;
  assign n5350 = n5349 ^ n5348;
  assign n5351 = ~n5222 & ~n5341;
  assign n5352 = ~n5346 & ~n5351;
  assign n5353 = n5352 ^ n5348;
  assign n5354 = ~n5350 & ~n5353;
  assign n5355 = n5354 ^ n5348;
  assign n5356 = ~n5343 & n5355;
  assign n5321 = n2449 & ~n3833;
  assign n5322 = n2459 & ~n3691;
  assign n5323 = ~n5321 & ~n5322;
  assign n5324 = n5323 ^ n595;
  assign n5325 = n1108 & n4066;
  assign n5326 = n5325 ^ n595;
  assign n5327 = n4066 & n4303;
  assign n5328 = n5327 ^ n595;
  assign n5329 = n595 & ~n5328;
  assign n5330 = n5329 ^ n595;
  assign n5331 = n5326 & n5330;
  assign n5332 = n5331 ^ n5329;
  assign n5333 = n5332 ^ n595;
  assign n5334 = n5333 ^ n5327;
  assign n5335 = ~n5324 & ~n5334;
  assign n5336 = n5335 ^ n5327;
  assign n5317 = n5255 ^ n5226;
  assign n5318 = n5233 & ~n5317;
  assign n5319 = n5318 ^ n5232;
  assign n5309 = n2320 ^ n812;
  assign n5310 = ~n5224 & n5309;
  assign n5311 = n5310 ^ n812;
  assign n5312 = n3150 & n5311;
  assign n5313 = ~n565 & ~n5312;
  assign n5314 = ~n3150 & ~n5311;
  assign n5315 = n5313 & ~n5314;
  assign n5295 = n596 & ~n4047;
  assign n5296 = ~n2488 & ~n3116;
  assign n5297 = n2492 & ~n3097;
  assign n5298 = ~n5296 & ~n5297;
  assign n5299 = ~n565 & n5298;
  assign n5300 = ~n5295 & n5299;
  assign n5301 = n4519 & n4596;
  assign n5302 = n3643 ^ n572;
  assign n5303 = n596 & ~n5302;
  assign n5304 = n3655 & n5303;
  assign n5305 = n565 & ~n5298;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = ~n5301 & n5306;
  assign n5308 = ~n5300 & n5307;
  assign n5316 = n5315 ^ n5308;
  assign n5320 = n5319 ^ n5316;
  assign n5337 = n5336 ^ n5320;
  assign n5357 = n5356 ^ n5337;
  assign n5286 = n866 & n3685;
  assign n5287 = n56 & ~n336;
  assign n5288 = n59 & ~n101;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n537 & n5289;
  assign n5291 = n883 & n928;
  assign n5292 = n5290 & n5291;
  assign n5293 = n5286 & n5292;
  assign n5294 = n396 & n5293;
  assign n5358 = n5357 ^ n5294;
  assign n5362 = n5361 ^ n5358;
  assign n5282 = n5183 & n5280;
  assign n5283 = ~n3797 & ~n5282;
  assign n5284 = n5194 & ~n5280;
  assign n5285 = ~n5283 & ~n5284;
  assign n5363 = n5362 ^ n5285;
  assign n5454 = n5361 ^ n5357;
  assign n5455 = ~n5358 & ~n5454;
  assign n5456 = n5455 ^ n5361;
  assign n5437 = n3814 ^ n595;
  assign n5438 = n5437 ^ n595;
  assign n5439 = ~n618 & ~n3833;
  assign n5440 = n5439 ^ n595;
  assign n5441 = ~n5438 & ~n5440;
  assign n5442 = n5441 ^ n595;
  assign n5443 = ~n2452 & ~n5442;
  assign n5444 = n2453 ^ n595;
  assign n5445 = n2453 ^ n618;
  assign n5446 = ~n5444 & n5445;
  assign n5447 = ~n3833 & n5446;
  assign n5448 = n5447 ^ n595;
  assign n5449 = ~n5443 & n5448;
  assign n5423 = n596 & ~n4707;
  assign n5424 = ~n2488 & n3643;
  assign n5425 = n2492 & ~n3116;
  assign n5426 = ~n5424 & ~n5425;
  assign n5427 = ~n565 & n5426;
  assign n5428 = ~n5423 & n5427;
  assign n5429 = n4261 & n4596;
  assign n5430 = n3691 ^ n572;
  assign n5431 = n596 & n5430;
  assign n5432 = n3676 & n5431;
  assign n5433 = n565 & ~n5426;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = ~n5429 & n5434;
  assign n5436 = ~n5428 & n5435;
  assign n5450 = n5449 ^ n5436;
  assign n5408 = ~n5219 & n5222;
  assign n5409 = ~n5338 & n5408;
  assign n5410 = ~n5337 & ~n5409;
  assign n5411 = ~n5205 & ~n5410;
  assign n5412 = n5219 & ~n5222;
  assign n5413 = n5337 & ~n5412;
  assign n5414 = ~n5340 & ~n5413;
  assign n5415 = ~n5411 & n5414;
  assign n5416 = n5337 & ~n5338;
  assign n5417 = n5222 ^ n5205;
  assign n5418 = n5219 ^ n5205;
  assign n5419 = ~n5417 & n5418;
  assign n5420 = n5419 ^ n5205;
  assign n5421 = ~n5416 & n5420;
  assign n5422 = ~n5415 & ~n5421;
  assign n5451 = n5450 ^ n5422;
  assign n5380 = ~n5308 & n5314;
  assign n5381 = ~n3097 & ~n5380;
  assign n5382 = n5308 & n5311;
  assign n5383 = n5248 & n5382;
  assign n5384 = n5381 & ~n5383;
  assign n5385 = n5313 & ~n5380;
  assign n5386 = n3150 & ~n5308;
  assign n5387 = n3097 & ~n5386;
  assign n5388 = ~n5385 & n5387;
  assign n5389 = ~n5384 & ~n5388;
  assign n5390 = n565 & ~n5308;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = n5336 ^ n5316;
  assign n5393 = ~n5320 & ~n5392;
  assign n5394 = n5393 ^ n5319;
  assign n5395 = ~n5391 & n5394;
  assign n5396 = ~n565 & ~n5314;
  assign n5397 = ~n5382 & n5396;
  assign n5398 = ~n5248 & n5308;
  assign n5399 = ~n3097 & ~n5398;
  assign n5400 = ~n5397 & n5399;
  assign n5401 = ~n565 & n5380;
  assign n5402 = n5308 & ~n5313;
  assign n5403 = n3097 & ~n5402;
  assign n5404 = ~n5401 & n5403;
  assign n5405 = ~n5400 & ~n5404;
  assign n5406 = ~n5394 & n5405;
  assign n5407 = ~n5395 & ~n5406;
  assign n5452 = n5451 ^ n5407;
  assign n5368 = ~n385 & ~n861;
  assign n5369 = ~n235 & ~n271;
  assign n5370 = ~n491 & n5369;
  assign n5371 = ~n5368 & n5370;
  assign n5372 = n109 & ~n123;
  assign n5373 = ~n205 & ~n5372;
  assign n5374 = n2111 & n5373;
  assign n5375 = n889 & n5374;
  assign n5376 = n4018 & n5375;
  assign n5377 = n1984 & n5376;
  assign n5378 = n194 & n5377;
  assign n5379 = n5371 & n5378;
  assign n5453 = n5452 ^ n5379;
  assign n5457 = n5456 ^ n5453;
  assign n5364 = n5282 & n5362;
  assign n5365 = ~n3797 & ~n5364;
  assign n5366 = n5284 & ~n5362;
  assign n5367 = ~n5365 & ~n5366;
  assign n5458 = n5457 ^ n5367;
  assign n5549 = n5456 ^ n5452;
  assign n5550 = n5453 & n5549;
  assign n5551 = n5550 ^ n5456;
  assign n5532 = n213 & n3469;
  assign n5533 = ~n363 & ~n465;
  assign n5534 = ~n319 & ~n2151;
  assign n5535 = n5533 & n5534;
  assign n5536 = n5532 & n5535;
  assign n5537 = ~n236 & ~n819;
  assign n5538 = n106 & ~n306;
  assign n5539 = ~n905 & ~n5538;
  assign n5540 = ~n5537 & n5539;
  assign n5541 = ~n197 & ~n214;
  assign n5542 = ~n3108 & n5541;
  assign n5543 = n5540 & n5542;
  assign n5544 = n5536 & n5543;
  assign n5545 = n833 & n5544;
  assign n5546 = n3432 & n5545;
  assign n5547 = n3967 & n5546;
  assign n5463 = ~n5395 & ~n5422;
  assign n5464 = ~n5406 & n5463;
  assign n5493 = ~n3097 & ~n3116;
  assign n5494 = n3097 & n3114;
  assign n5495 = ~n565 & ~n5494;
  assign n5496 = ~n5493 & n5495;
  assign n5497 = n5496 ^ n595;
  assign n5467 = n3833 ^ n572;
  assign n5468 = n3815 & n5467;
  assign n5469 = ~n4381 & ~n5468;
  assign n5470 = n2301 & n3643;
  assign n5471 = ~n2488 & ~n3691;
  assign n5472 = ~n565 & ~n5471;
  assign n5473 = ~n5470 & n5472;
  assign n5474 = ~n5469 & n5473;
  assign n5475 = n3691 ^ n565;
  assign n5476 = n611 & n5475;
  assign n5477 = ~n572 & ~n5476;
  assign n5478 = n2490 & ~n3643;
  assign n5479 = n5478 ^ n2478;
  assign n5480 = n5477 & ~n5479;
  assign n5481 = n2475 & ~n3643;
  assign n5482 = n2490 & ~n3691;
  assign n5483 = n572 & ~n5482;
  assign n5484 = ~n5481 & n5483;
  assign n5485 = ~n5480 & ~n5484;
  assign n5486 = ~n565 & n3691;
  assign n5487 = n2478 & n5486;
  assign n5488 = ~n5485 & ~n5487;
  assign n5489 = ~n5474 & n5488;
  assign n5490 = ~n4393 & ~n5468;
  assign n5491 = n4596 & ~n5490;
  assign n5492 = n5489 & ~n5491;
  assign n5498 = n5497 ^ n5492;
  assign n5465 = ~n565 & n5381;
  assign n5466 = ~n5402 & ~n5465;
  assign n5499 = n5498 ^ n5466;
  assign n5500 = ~n5406 & ~n5499;
  assign n5501 = n5422 & ~n5500;
  assign n5502 = ~n5464 & ~n5501;
  assign n5503 = ~n5395 & n5499;
  assign n5504 = ~n5436 & n5449;
  assign n5505 = ~n5503 & ~n5504;
  assign n5506 = ~n5502 & n5505;
  assign n5507 = ~n5422 & ~n5499;
  assign n5508 = n5499 ^ n5406;
  assign n5509 = n5436 & ~n5449;
  assign n5510 = n5509 ^ n5504;
  assign n5511 = n5510 ^ n5504;
  assign n5512 = n5504 ^ n5499;
  assign n5513 = n5512 ^ n5504;
  assign n5514 = n5511 & n5513;
  assign n5515 = n5514 ^ n5504;
  assign n5516 = n5508 & n5515;
  assign n5517 = n5516 ^ n5504;
  assign n5518 = ~n5507 & n5517;
  assign n5519 = ~n5464 & n5518;
  assign n5520 = n5463 & ~n5499;
  assign n5521 = n5509 & n5520;
  assign n5522 = ~n5519 & ~n5521;
  assign n5523 = ~n5506 & n5522;
  assign n5524 = n5463 & n5504;
  assign n5525 = ~n5407 & n5422;
  assign n5526 = ~n5406 & n5499;
  assign n5527 = ~n5509 & ~n5526;
  assign n5528 = ~n5525 & n5527;
  assign n5529 = ~n5524 & ~n5528;
  assign n5530 = ~n5520 & ~n5529;
  assign n5531 = n5523 & ~n5530;
  assign n5548 = n5547 ^ n5531;
  assign n5552 = n5551 ^ n5548;
  assign n5459 = n5364 & ~n5457;
  assign n5460 = ~n3797 & ~n5459;
  assign n5461 = n5366 & n5457;
  assign n5462 = ~n5460 & ~n5461;
  assign n5553 = n5552 ^ n5462;
  assign n5604 = n5551 ^ n5531;
  assign n5605 = ~n5548 & ~n5604;
  assign n5606 = n5605 ^ n5551;
  assign n5591 = ~n267 & ~n399;
  assign n5592 = n2111 & n5591;
  assign n5593 = n86 & ~n5039;
  assign n5594 = n5592 & ~n5593;
  assign n5595 = ~n173 & ~n1964;
  assign n5596 = n361 & n5595;
  assign n5597 = n3106 & n5596;
  assign n5598 = n5594 & n5597;
  assign n5599 = n896 & n5598;
  assign n5600 = n1287 & n5599;
  assign n5601 = n1915 & n2292;
  assign n5602 = n5600 & n5601;
  assign n5586 = n5492 ^ n5466;
  assign n5587 = ~n5498 & ~n5586;
  assign n5588 = n5587 ^ n5466;
  assign n5581 = ~n595 & ~n5494;
  assign n5582 = ~n5493 & ~n5581;
  assign n5583 = n5582 ^ n3643;
  assign n5584 = ~n565 & n5583;
  assign n5567 = n573 & n4066;
  assign n5568 = n596 & ~n5567;
  assign n5569 = n572 & ~n3833;
  assign n5570 = n2507 & ~n3691;
  assign n5571 = n2478 & ~n5570;
  assign n5572 = ~n5569 & n5571;
  assign n5573 = n5467 ^ n3833;
  assign n5574 = ~n565 & ~n3691;
  assign n5575 = n5574 ^ n3833;
  assign n5576 = n5573 & ~n5575;
  assign n5577 = n5576 ^ n3833;
  assign n5578 = n611 & n5577;
  assign n5579 = ~n5572 & ~n5578;
  assign n5580 = ~n5568 & n5579;
  assign n5585 = n5584 ^ n5580;
  assign n5589 = n5588 ^ n5585;
  assign n5558 = ~n5503 & n5509;
  assign n5559 = ~n5500 & ~n5558;
  assign n5560 = ~n5422 & n5559;
  assign n5561 = n5503 & ~n5509;
  assign n5562 = n5508 & ~n5512;
  assign n5563 = n5562 ^ n5406;
  assign n5564 = ~n5561 & ~n5563;
  assign n5565 = ~n5560 & n5564;
  assign n5566 = ~n5524 & n5565;
  assign n5590 = n5589 ^ n5566;
  assign n5603 = n5602 ^ n5590;
  assign n5607 = n5606 ^ n5603;
  assign n5554 = n5459 & n5552;
  assign n5555 = ~n3797 & ~n5554;
  assign n5556 = n5461 & ~n5552;
  assign n5557 = ~n5555 & ~n5556;
  assign n5608 = n5607 ^ n5557;
  assign n5683 = n5606 ^ n5590;
  assign n5684 = n5603 & n5683;
  assign n5685 = n5684 ^ n5606;
  assign n5626 = n5588 ^ n5566;
  assign n5627 = n5589 & ~n5626;
  assign n5628 = n5627 ^ n5566;
  assign n5642 = n3643 & n5574;
  assign n5643 = n5580 ^ n3643;
  assign n5644 = n5583 & n5643;
  assign n5645 = n5644 ^ n3643;
  assign n5646 = ~n565 & ~n5645;
  assign n5647 = n5642 & n5646;
  assign n5637 = n5580 & n5582;
  assign n5629 = n596 & n3814;
  assign n5630 = n573 & n2488;
  assign n5631 = ~n3833 & n5630;
  assign n5632 = ~n5629 & n5631;
  assign n5633 = ~n3643 & ~n5632;
  assign n5666 = n5486 & n5633;
  assign n5667 = ~n5637 & n5666;
  assign n5668 = ~n5647 & ~n5667;
  assign n5648 = ~n3643 & n3691;
  assign n5669 = n5632 & ~n5648;
  assign n5654 = n5645 ^ n5580;
  assign n5655 = ~n565 & ~n5654;
  assign n5656 = n5655 ^ n5580;
  assign n5670 = n5669 ^ n5656;
  assign n5671 = n5670 ^ n5669;
  assign n5672 = n3691 ^ n3643;
  assign n5673 = ~n565 & n5672;
  assign n5674 = ~n5632 & ~n5673;
  assign n5675 = n5674 ^ n5669;
  assign n5676 = ~n5671 & n5675;
  assign n5677 = n5676 ^ n5669;
  assign n5678 = n5668 & ~n5677;
  assign n5634 = ~n3691 & n5633;
  assign n5635 = n5580 ^ n565;
  assign n5636 = n5635 ^ n5580;
  assign n5638 = n5637 ^ n5580;
  assign n5639 = ~n5636 & ~n5638;
  assign n5640 = n5639 ^ n5580;
  assign n5641 = n5634 & n5640;
  assign n5649 = n565 & ~n5580;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = ~n5647 & n5650;
  assign n5652 = n5651 ^ n5632;
  assign n5653 = n5652 ^ n5651;
  assign n5657 = ~n565 & ~n3643;
  assign n5658 = ~n5574 & ~n5657;
  assign n5659 = n5656 & n5658;
  assign n5660 = n5642 & ~n5646;
  assign n5661 = ~n5659 & ~n5660;
  assign n5662 = n5661 ^ n5651;
  assign n5663 = ~n5653 & n5662;
  assign n5664 = n5663 ^ n5651;
  assign n5665 = ~n5641 & n5664;
  assign n5679 = n5678 ^ n5665;
  assign n5680 = ~n5628 & n5679;
  assign n5681 = n5680 ^ n5665;
  assign n5613 = ~n472 & n897;
  assign n5614 = n1062 & n5613;
  assign n5615 = ~n93 & ~n647;
  assign n5616 = n5595 & n5615;
  assign n5617 = n60 & ~n454;
  assign n5618 = ~n426 & ~n5617;
  assign n5619 = ~n923 & n5618;
  assign n5620 = n5616 & n5619;
  assign n5621 = n3440 & n5620;
  assign n5622 = n1011 & n5621;
  assign n5623 = n2118 & n5622;
  assign n5624 = n5614 & n5623;
  assign n5625 = n5371 & n5624;
  assign n5682 = n5681 ^ n5625;
  assign n5686 = n5685 ^ n5682;
  assign n5609 = n5556 & n5607;
  assign n5610 = n3797 & ~n5609;
  assign n5611 = n5554 & ~n5607;
  assign n5612 = ~n5610 & ~n5611;
  assign n5687 = n5686 ^ n5612;
  assign n5725 = n5685 ^ n5681;
  assign n5726 = n5682 & n5725;
  assign n5727 = n5726 ^ n5685;
  assign n5713 = ~n60 & n1985;
  assign n5714 = ~n2146 & ~n5713;
  assign n5715 = ~n438 & ~n1964;
  assign n5716 = ~n521 & n5715;
  assign n5717 = n3431 & n5716;
  assign n5718 = n3082 & n5717;
  assign n5719 = n3511 & n5718;
  assign n5720 = n5535 & n5719;
  assign n5721 = n3445 & n5720;
  assign n5722 = n877 & n5721;
  assign n5723 = ~n5714 & n5722;
  assign n5705 = n565 & ~n5632;
  assign n5706 = n572 & n3691;
  assign n5707 = n5481 & n5706;
  assign n5708 = n3643 & ~n5486;
  assign n5709 = n3833 & ~n5708;
  assign n5710 = ~n5707 & ~n5709;
  assign n5711 = ~n5705 & n5710;
  assign n5692 = n3691 & n5632;
  assign n5693 = n5692 ^ n5673;
  assign n5694 = n5692 ^ n5656;
  assign n5695 = ~n5692 & ~n5694;
  assign n5696 = n5695 ^ n5692;
  assign n5697 = ~n5693 & ~n5696;
  assign n5698 = n5697 ^ n5695;
  assign n5699 = n5698 ^ n5692;
  assign n5700 = n5699 ^ n5656;
  assign n5701 = ~n5669 & ~n5700;
  assign n5702 = n5628 & ~n5701;
  assign n5703 = ~n5656 & ~n5674;
  assign n5704 = ~n5702 & ~n5703;
  assign n5712 = n5711 ^ n5704;
  assign n5724 = n5723 ^ n5712;
  assign n5728 = n5727 ^ n5724;
  assign n5688 = n5611 & ~n5686;
  assign n5689 = ~n3797 & ~n5688;
  assign n5690 = n5609 & n5686;
  assign n5691 = ~n5689 & ~n5690;
  assign n5729 = n5728 ^ n5691;
  assign n5745 = n5727 ^ n5712;
  assign n5746 = ~n5724 & ~n5745;
  assign n5747 = n5746 ^ n5727;
  assign n5734 = n714 & n1932;
  assign n5735 = n5541 & n5734;
  assign n5736 = ~n174 & ~n727;
  assign n5737 = n276 & n5736;
  assign n5738 = n196 & ~n219;
  assign n5739 = ~n385 & ~n5738;
  assign n5740 = n872 & ~n5739;
  assign n5741 = n5737 & n5740;
  assign n5742 = n5735 & n5741;
  assign n5743 = n531 & n5742;
  assign n5744 = n3093 & n5743;
  assign n5748 = n5747 ^ n5744;
  assign n5730 = n5690 & ~n5728;
  assign n5731 = n3797 & ~n5730;
  assign n5732 = n5688 & n5728;
  assign n5733 = ~n5731 & ~n5732;
  assign n5749 = n5748 ^ n5733;
  assign n5760 = n822 & n908;
  assign n5761 = n370 & ~n931;
  assign n5762 = n3509 & n4337;
  assign n5763 = n5761 & n5762;
  assign n5764 = n1068 & n5763;
  assign n5765 = n5760 & n5764;
  assign n5766 = n487 & n5765;
  assign n5767 = n1003 & n5766;
  assign n5768 = n3459 & n5767;
  assign n5750 = n5747 ^ n5732;
  assign n5751 = n5748 & n5750;
  assign n5752 = n5751 ^ n5732;
  assign n5753 = ~n3797 & ~n5752;
  assign n5754 = n5744 & ~n5747;
  assign n5755 = n5730 & n5754;
  assign n5756 = ~n5744 & n5747;
  assign n5757 = n5731 & n5756;
  assign n5758 = ~n5755 & ~n5757;
  assign n5759 = ~n5753 & n5758;
  assign n5769 = n5768 ^ n5759;
  assign n5778 = n106 & ~n3085;
  assign n5779 = n188 & ~n5778;
  assign n5780 = n110 & n335;
  assign n5781 = ~n371 & ~n5780;
  assign n5782 = n5779 & n5781;
  assign n5783 = n4624 & n5782;
  assign n5784 = n2392 & n5783;
  assign n5785 = n859 & n5784;
  assign n5786 = n5614 & n5785;
  assign n5777 = n5752 & ~n5768;
  assign n5787 = n5786 ^ n5777;
  assign n5770 = ~n5756 & ~n5768;
  assign n5771 = n5730 & ~n5770;
  assign n5772 = n5732 & ~n5748;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = ~n5755 & n5768;
  assign n5775 = ~n5773 & ~n5774;
  assign n5776 = n3797 & ~n5775;
  assign n5788 = n5787 ^ n5776;
  assign n5799 = n5786 ^ n5775;
  assign n5800 = n5799 ^ n5786;
  assign n5801 = n5786 ^ n3797;
  assign n5802 = n5801 ^ n5786;
  assign n5803 = n5800 & n5802;
  assign n5804 = n5803 ^ n5786;
  assign n5805 = n5787 & ~n5804;
  assign n5806 = n5805 ^ n3797;
  assign n5789 = ~n172 & ~n501;
  assign n5790 = ~n204 & n5789;
  assign n5791 = ~n444 & n5790;
  assign n5792 = n163 & n904;
  assign n5793 = ~n225 & ~n5792;
  assign n5794 = n5791 & ~n5793;
  assign n5795 = n4631 & n5794;
  assign n5796 = ~n3101 & n5795;
  assign n5797 = n912 & n5796;
  assign n5798 = n5043 & n5797;
  assign n5807 = n5806 ^ n5798;
  assign n5814 = n5777 ^ n3797;
  assign n5815 = ~n5786 & ~n5798;
  assign n5816 = n5815 ^ n5777;
  assign n5817 = n5816 ^ n5815;
  assign n5818 = n5786 & n5798;
  assign n5819 = n5818 ^ n5815;
  assign n5820 = ~n5817 & n5819;
  assign n5821 = n5820 ^ n5815;
  assign n5822 = n5814 & n5821;
  assign n5823 = n5822 ^ n3797;
  assign n5824 = n5823 ^ n5798;
  assign n5825 = n5824 ^ n5823;
  assign n5826 = n5777 & ~n5786;
  assign n5827 = n5826 ^ n5823;
  assign n5828 = n5827 ^ n5823;
  assign n5829 = ~n5825 & n5828;
  assign n5830 = n5829 ^ n5823;
  assign n5831 = n5776 & ~n5830;
  assign n5832 = n5831 ^ n5823;
  assign n5808 = ~n59 & n115;
  assign n5809 = ~n532 & ~n5808;
  assign n5810 = ~n459 & ~n473;
  assign n5811 = n318 & n5810;
  assign n5812 = n3631 & n5811;
  assign n5813 = ~n5809 & n5812;
  assign n5833 = n5832 ^ n5813;
  assign n5835 = ~n5813 & n5815;
  assign n5836 = n5777 & n5835;
  assign n5834 = n804 & ~n3638;
  assign n5840 = n5836 ^ n5834;
  assign n5841 = n5840 ^ n3797;
  assign n5837 = n5836 ^ n5777;
  assign n5838 = ~n5834 & ~n5837;
  assign n5839 = n5838 ^ n5777;
  assign n5842 = n5841 ^ n5839;
  assign n5843 = n5840 ^ n5839;
  assign n5844 = n5813 & n5818;
  assign n5845 = n5844 ^ n5835;
  assign n5846 = ~n5777 & n5845;
  assign n5847 = n5846 ^ n5835;
  assign n5848 = n5775 & n5847;
  assign n5849 = n5848 ^ n5840;
  assign n5850 = ~n5840 & ~n5849;
  assign n5851 = n5850 ^ n5840;
  assign n5852 = n5843 & ~n5851;
  assign n5853 = n5852 ^ n5850;
  assign n5854 = n5853 ^ n5840;
  assign n5855 = n5854 ^ n5848;
  assign n5856 = ~n5842 & ~n5855;
  assign n5857 = n5856 ^ n5841;
  assign n5858 = ~x21 & ~x22;
  assign n5859 = n804 & n5858;
  assign n5860 = ~n5834 & n5836;
  assign n5861 = n5776 ^ n3797;
  assign n5862 = n5860 & ~n5861;
  assign n5863 = n5862 ^ n3797;
  assign n5864 = ~n5859 & ~n5863;
  assign n5865 = n5834 & ~n5836;
  assign n5866 = ~n5858 & n5865;
  assign n5867 = n5848 & n5866;
  assign n5868 = ~n5864 & ~n5867;
  assign n5869 = n3797 & ~n5867;
  assign y0 = ~n3796;
  assign y1 = n3970;
  assign y2 = ~n4164;
  assign y3 = ~n4349;
  assign y4 = n4479;
  assign y5 = n4656;
  assign y6 = n4797;
  assign y7 = n4917;
  assign y8 = ~n5057;
  assign y9 = ~n5174;
  assign y10 = n5281;
  assign y11 = n5363;
  assign y12 = ~n5458;
  assign y13 = n5553;
  assign y14 = ~n5608;
  assign y15 = n5687;
  assign y16 = n5729;
  assign y17 = n5749;
  assign y18 = ~n5769;
  assign y19 = ~n5788;
  assign y20 = ~n5807;
  assign y21 = ~n5833;
  assign y22 = ~n5857;
  assign y23 = n5868;
  assign y24 = n5869;
endmodule