module Xor(
    //output logic out
);

    logic a;
    logic b;

    assign a = 0;
    assign b = a;

    //assign out = a ^ b;
    
endmodule
