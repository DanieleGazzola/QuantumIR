module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922;
  assign n514 = x383 & x511;
  assign n513 = x127 & x255;
  assign n515 = n514 ^ n513;
  assign n1063 = x510 ^ x382;
  assign n1064 = x511 ^ x383;
  assign n1065 = x509 ^ x381;
  assign n1066 = x380 & ~x508;
  assign n1067 = n1066 ^ x509;
  assign n1068 = ~n1065 & ~n1067;
  assign n1069 = n1068 ^ x509;
  assign n1070 = n1069 ^ x510;
  assign n1071 = ~n1063 & n1070;
  assign n1072 = n1071 ^ x510;
  assign n1073 = n1072 ^ x511;
  assign n1074 = n1073 ^ x511;
  assign n1075 = ~x381 & x509;
  assign n1076 = ~x382 & x510;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~x379 & x507;
  assign n1079 = ~x380 & x508;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = n1077 & n1080;
  assign n1082 = x379 & ~x507;
  assign n1083 = x506 ^ x378;
  assign n1084 = x505 ^ x377;
  assign n1085 = x504 ^ x376;
  assign n1086 = x503 ^ x375;
  assign n1087 = x502 ^ x374;
  assign n1088 = x501 ^ x373;
  assign n1089 = x500 ^ x372;
  assign n1090 = x499 ^ x371;
  assign n1091 = x498 ^ x370;
  assign n1092 = x497 ^ x369;
  assign n1093 = x496 ^ x368;
  assign n1094 = x495 ^ x367;
  assign n1095 = x494 ^ x366;
  assign n1096 = x493 ^ x365;
  assign n1097 = x492 ^ x364;
  assign n1098 = x491 ^ x363;
  assign n1099 = x490 ^ x362;
  assign n1100 = x489 ^ x361;
  assign n1101 = x488 ^ x360;
  assign n1102 = x487 ^ x359;
  assign n1103 = x486 ^ x358;
  assign n1104 = x485 ^ x357;
  assign n1105 = x484 ^ x356;
  assign n1106 = x483 ^ x355;
  assign n1107 = x482 ^ x354;
  assign n1108 = x481 ^ x353;
  assign n1109 = x480 ^ x352;
  assign n1110 = x479 ^ x351;
  assign n1111 = x478 ^ x350;
  assign n1112 = x477 ^ x349;
  assign n1113 = x476 ^ x348;
  assign n1114 = x475 ^ x347;
  assign n1115 = x474 ^ x346;
  assign n1116 = x473 ^ x345;
  assign n1117 = x472 ^ x344;
  assign n1118 = x471 ^ x343;
  assign n1119 = x470 ^ x342;
  assign n1120 = x469 ^ x341;
  assign n1121 = x468 ^ x340;
  assign n1122 = x467 ^ x339;
  assign n1123 = x466 ^ x338;
  assign n1124 = x465 ^ x337;
  assign n1125 = x464 ^ x336;
  assign n1126 = x463 ^ x335;
  assign n1127 = x462 ^ x334;
  assign n1128 = x461 ^ x333;
  assign n1129 = x460 ^ x332;
  assign n1130 = x459 ^ x331;
  assign n1131 = x458 ^ x330;
  assign n1132 = x457 ^ x329;
  assign n1133 = x456 ^ x328;
  assign n1134 = ~x327 & x455;
  assign n1135 = n1134 ^ x456;
  assign n1136 = n1135 ^ x456;
  assign n1137 = ~x325 & x453;
  assign n1138 = ~x326 & x454;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~x323 & x451;
  assign n1141 = ~x324 & x452;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = n1139 & n1142;
  assign n1144 = x323 & ~x451;
  assign n1145 = x450 ^ x322;
  assign n1146 = x449 ^ x321;
  assign n1147 = ~x320 & x448;
  assign n1148 = n1147 ^ x449;
  assign n1149 = n1148 ^ x449;
  assign n1150 = x315 & ~x443;
  assign n1151 = x442 ^ x314;
  assign n1152 = x441 ^ x313;
  assign n1153 = x440 ^ x312;
  assign n1154 = x439 ^ x311;
  assign n1155 = x438 ^ x310;
  assign n1156 = x437 ^ x309;
  assign n1157 = x436 ^ x308;
  assign n1158 = ~x307 & x435;
  assign n1159 = n1158 ^ x436;
  assign n1160 = n1159 ^ x436;
  assign n1161 = ~x297 & x425;
  assign n1162 = ~x298 & x426;
  assign n1163 = ~n1161 & ~n1162;
  assign n1164 = ~x295 & x423;
  assign n1165 = ~x296 & x424;
  assign n1166 = ~n1164 & ~n1165;
  assign n1167 = n1163 & n1166;
  assign n1168 = x295 & ~x423;
  assign n1169 = x422 ^ x294;
  assign n1170 = x421 ^ x293;
  assign n1171 = x420 ^ x292;
  assign n1172 = x419 ^ x291;
  assign n1173 = x418 ^ x290;
  assign n1174 = x417 ^ x289;
  assign n1175 = x416 ^ x288;
  assign n1176 = x415 ^ x287;
  assign n1177 = x414 ^ x286;
  assign n1178 = x413 ^ x285;
  assign n1179 = x412 ^ x284;
  assign n1180 = x411 ^ x283;
  assign n1181 = x410 ^ x282;
  assign n1182 = x409 ^ x281;
  assign n1183 = x408 ^ x280;
  assign n1184 = x407 ^ x279;
  assign n1185 = x406 ^ x278;
  assign n1186 = x405 ^ x277;
  assign n1187 = x404 ^ x276;
  assign n1188 = x403 ^ x275;
  assign n1189 = x402 ^ x274;
  assign n1190 = x401 ^ x273;
  assign n1191 = x400 ^ x272;
  assign n1192 = x399 ^ x271;
  assign n1193 = x398 ^ x270;
  assign n1194 = x397 ^ x269;
  assign n1195 = x396 ^ x268;
  assign n1196 = x395 ^ x267;
  assign n1197 = x394 ^ x266;
  assign n1198 = x393 ^ x265;
  assign n1199 = x392 ^ x264;
  assign n1200 = x391 ^ x263;
  assign n1201 = x390 ^ x262;
  assign n1202 = x389 ^ x261;
  assign n1203 = x388 ^ x260;
  assign n1204 = x387 ^ x259;
  assign n1205 = x386 ^ x258;
  assign n1206 = x385 ^ x257;
  assign n1207 = x256 & ~x384;
  assign n1208 = n1207 ^ x385;
  assign n1209 = ~n1206 & ~n1208;
  assign n1210 = n1209 ^ x385;
  assign n1211 = n1210 ^ x386;
  assign n1212 = ~n1205 & n1211;
  assign n1213 = n1212 ^ x386;
  assign n1214 = n1213 ^ x387;
  assign n1215 = ~n1204 & ~n1214;
  assign n1216 = n1215 ^ x259;
  assign n1217 = n1216 ^ x388;
  assign n1218 = ~n1203 & n1217;
  assign n1219 = n1218 ^ x260;
  assign n1220 = n1219 ^ x389;
  assign n1221 = ~n1202 & ~n1220;
  assign n1222 = n1221 ^ x389;
  assign n1223 = n1222 ^ x390;
  assign n1224 = ~n1201 & n1223;
  assign n1225 = n1224 ^ x390;
  assign n1226 = n1225 ^ x391;
  assign n1227 = ~n1200 & n1226;
  assign n1228 = n1227 ^ x391;
  assign n1229 = n1228 ^ x392;
  assign n1230 = ~n1199 & n1229;
  assign n1231 = n1230 ^ x392;
  assign n1232 = n1231 ^ x393;
  assign n1233 = ~n1198 & n1232;
  assign n1234 = n1233 ^ x393;
  assign n1235 = n1234 ^ x394;
  assign n1236 = ~n1197 & ~n1235;
  assign n1237 = n1236 ^ x266;
  assign n1238 = n1237 ^ x395;
  assign n1239 = ~n1196 & n1238;
  assign n1240 = n1239 ^ x267;
  assign n1241 = n1240 ^ x396;
  assign n1242 = ~n1195 & n1241;
  assign n1243 = n1242 ^ x268;
  assign n1244 = n1243 ^ x397;
  assign n1245 = ~n1194 & n1244;
  assign n1246 = n1245 ^ x269;
  assign n1247 = n1246 ^ x398;
  assign n1248 = ~n1193 & n1247;
  assign n1249 = n1248 ^ x270;
  assign n1250 = n1249 ^ x399;
  assign n1251 = ~n1192 & n1250;
  assign n1252 = n1251 ^ x271;
  assign n1253 = n1252 ^ x400;
  assign n1254 = ~n1191 & n1253;
  assign n1255 = n1254 ^ x272;
  assign n1256 = n1255 ^ x401;
  assign n1257 = ~n1190 & n1256;
  assign n1258 = n1257 ^ x273;
  assign n1259 = n1258 ^ x402;
  assign n1260 = ~n1189 & ~n1259;
  assign n1261 = n1260 ^ x402;
  assign n1262 = n1261 ^ x403;
  assign n1263 = ~n1188 & ~n1262;
  assign n1264 = n1263 ^ x275;
  assign n1265 = n1264 ^ x404;
  assign n1266 = ~n1187 & n1265;
  assign n1267 = n1266 ^ x276;
  assign n1268 = n1267 ^ x405;
  assign n1269 = ~n1186 & ~n1268;
  assign n1270 = n1269 ^ x405;
  assign n1271 = n1270 ^ x406;
  assign n1272 = ~n1185 & n1271;
  assign n1273 = n1272 ^ x406;
  assign n1274 = n1273 ^ x407;
  assign n1275 = ~n1184 & n1274;
  assign n1276 = n1275 ^ x407;
  assign n1277 = n1276 ^ x408;
  assign n1278 = ~n1183 & n1277;
  assign n1279 = n1278 ^ x408;
  assign n1280 = n1279 ^ x409;
  assign n1281 = ~n1182 & ~n1280;
  assign n1282 = n1281 ^ x281;
  assign n1283 = n1282 ^ x410;
  assign n1284 = ~n1181 & n1283;
  assign n1285 = n1284 ^ x282;
  assign n1286 = n1285 ^ x411;
  assign n1287 = ~n1180 & ~n1286;
  assign n1288 = n1287 ^ x411;
  assign n1289 = n1288 ^ x412;
  assign n1290 = ~n1179 & n1289;
  assign n1291 = n1290 ^ x412;
  assign n1292 = n1291 ^ x413;
  assign n1293 = ~n1178 & ~n1292;
  assign n1294 = n1293 ^ x285;
  assign n1295 = n1294 ^ x414;
  assign n1296 = ~n1177 & n1295;
  assign n1297 = n1296 ^ x286;
  assign n1298 = n1297 ^ x415;
  assign n1299 = ~n1176 & ~n1298;
  assign n1300 = n1299 ^ x415;
  assign n1301 = n1300 ^ x416;
  assign n1302 = ~n1175 & n1301;
  assign n1303 = n1302 ^ x416;
  assign n1304 = n1303 ^ x417;
  assign n1305 = ~n1174 & n1304;
  assign n1306 = n1305 ^ x417;
  assign n1307 = n1306 ^ x418;
  assign n1308 = ~n1173 & ~n1307;
  assign n1309 = n1308 ^ x290;
  assign n1310 = n1309 ^ x419;
  assign n1311 = ~n1172 & n1310;
  assign n1312 = n1311 ^ x291;
  assign n1313 = n1312 ^ x420;
  assign n1314 = ~n1171 & n1313;
  assign n1315 = n1314 ^ x292;
  assign n1316 = n1315 ^ x421;
  assign n1317 = ~n1170 & n1316;
  assign n1318 = n1317 ^ x293;
  assign n1319 = n1318 ^ x422;
  assign n1320 = ~n1169 & ~n1319;
  assign n1321 = n1320 ^ x422;
  assign n1322 = ~n1168 & n1321;
  assign n1323 = n1167 & ~n1322;
  assign n1324 = x299 & ~x427;
  assign n1325 = x426 ^ x298;
  assign n1326 = x425 ^ x297;
  assign n1327 = x296 & ~x424;
  assign n1328 = n1327 ^ x425;
  assign n1329 = ~n1326 & ~n1328;
  assign n1330 = n1329 ^ x425;
  assign n1331 = n1330 ^ x426;
  assign n1332 = ~n1325 & n1331;
  assign n1333 = n1332 ^ x426;
  assign n1334 = ~n1324 & n1333;
  assign n1335 = ~n1323 & n1334;
  assign n1336 = ~x302 & x430;
  assign n1337 = ~x301 & x429;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~x299 & x427;
  assign n1340 = ~x300 & x428;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = n1338 & n1341;
  assign n1343 = ~n1335 & n1342;
  assign n1344 = x303 & ~x431;
  assign n1345 = x430 ^ x302;
  assign n1346 = x429 ^ x301;
  assign n1347 = x300 & ~x428;
  assign n1348 = n1347 ^ x429;
  assign n1349 = ~n1346 & ~n1348;
  assign n1350 = n1349 ^ x429;
  assign n1351 = n1350 ^ x430;
  assign n1352 = ~n1345 & n1351;
  assign n1353 = n1352 ^ x430;
  assign n1354 = ~n1344 & n1353;
  assign n1355 = ~n1343 & n1354;
  assign n1356 = ~x304 & x432;
  assign n1357 = ~x303 & x431;
  assign n1358 = ~n1356 & ~n1357;
  assign n1359 = ~n1355 & n1358;
  assign n1360 = x305 & ~x433;
  assign n1361 = x304 & ~x432;
  assign n1362 = ~n1360 & ~n1361;
  assign n1363 = ~n1359 & n1362;
  assign n1364 = ~x306 & x434;
  assign n1365 = ~x305 & x433;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1363 & n1366;
  assign n1368 = x307 & ~x435;
  assign n1369 = x306 & ~x434;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~n1367 & n1370;
  assign n1372 = n1371 ^ x436;
  assign n1373 = n1372 ^ x436;
  assign n1374 = ~n1160 & ~n1373;
  assign n1375 = n1374 ^ x436;
  assign n1376 = ~n1157 & n1375;
  assign n1377 = n1376 ^ x308;
  assign n1378 = n1377 ^ x437;
  assign n1379 = ~n1156 & ~n1378;
  assign n1380 = n1379 ^ x437;
  assign n1381 = n1380 ^ x438;
  assign n1382 = ~n1155 & n1381;
  assign n1383 = n1382 ^ x438;
  assign n1384 = n1383 ^ x439;
  assign n1385 = ~n1154 & n1384;
  assign n1386 = n1385 ^ x439;
  assign n1387 = n1386 ^ x440;
  assign n1388 = ~n1153 & n1387;
  assign n1389 = n1388 ^ x440;
  assign n1390 = n1389 ^ x441;
  assign n1391 = ~n1152 & ~n1390;
  assign n1392 = n1391 ^ x313;
  assign n1393 = n1392 ^ x442;
  assign n1394 = ~n1151 & n1393;
  assign n1395 = n1394 ^ x314;
  assign n1396 = ~n1150 & ~n1395;
  assign n1397 = ~x315 & x443;
  assign n1398 = ~x316 & x444;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~x318 & x446;
  assign n1401 = ~x317 & x445;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~x319 & x447;
  assign n1404 = n1402 & ~n1403;
  assign n1405 = n1399 & n1404;
  assign n1406 = ~n1396 & n1405;
  assign n1407 = x317 & ~x445;
  assign n1408 = x316 & ~x444;
  assign n1409 = ~n1407 & ~n1408;
  assign n1410 = n1404 & ~n1409;
  assign n1411 = x320 & ~x448;
  assign n1412 = x447 ^ x319;
  assign n1413 = x318 & ~x446;
  assign n1414 = n1413 ^ x447;
  assign n1415 = ~n1412 & n1414;
  assign n1416 = n1415 ^ x319;
  assign n1417 = ~n1411 & ~n1416;
  assign n1418 = ~n1410 & n1417;
  assign n1419 = ~n1406 & n1418;
  assign n1420 = n1419 ^ x449;
  assign n1421 = n1420 ^ x449;
  assign n1422 = ~n1149 & ~n1421;
  assign n1423 = n1422 ^ x449;
  assign n1424 = ~n1146 & n1423;
  assign n1425 = n1424 ^ x321;
  assign n1426 = n1425 ^ x450;
  assign n1427 = ~n1145 & ~n1426;
  assign n1428 = n1427 ^ x450;
  assign n1429 = ~n1144 & n1428;
  assign n1430 = n1143 & ~n1429;
  assign n1431 = x327 & ~x455;
  assign n1432 = x454 ^ x326;
  assign n1433 = x453 ^ x325;
  assign n1434 = x324 & ~x452;
  assign n1435 = n1434 ^ x453;
  assign n1436 = ~n1433 & ~n1435;
  assign n1437 = n1436 ^ x453;
  assign n1438 = n1437 ^ x454;
  assign n1439 = ~n1432 & n1438;
  assign n1440 = n1439 ^ x454;
  assign n1441 = ~n1431 & n1440;
  assign n1442 = ~n1430 & n1441;
  assign n1443 = n1442 ^ x456;
  assign n1444 = n1443 ^ x456;
  assign n1445 = ~n1136 & ~n1444;
  assign n1446 = n1445 ^ x456;
  assign n1447 = ~n1133 & n1446;
  assign n1448 = n1447 ^ x328;
  assign n1449 = n1448 ^ x457;
  assign n1450 = ~n1132 & ~n1449;
  assign n1451 = n1450 ^ x457;
  assign n1452 = n1451 ^ x458;
  assign n1453 = ~n1131 & ~n1452;
  assign n1454 = n1453 ^ x330;
  assign n1455 = n1454 ^ x459;
  assign n1456 = ~n1130 & n1455;
  assign n1457 = n1456 ^ x331;
  assign n1458 = n1457 ^ x460;
  assign n1459 = ~n1129 & ~n1458;
  assign n1460 = n1459 ^ x460;
  assign n1461 = n1460 ^ x461;
  assign n1462 = ~n1128 & ~n1461;
  assign n1463 = n1462 ^ x333;
  assign n1464 = n1463 ^ x462;
  assign n1465 = ~n1127 & n1464;
  assign n1466 = n1465 ^ x334;
  assign n1467 = n1466 ^ x463;
  assign n1468 = ~n1126 & ~n1467;
  assign n1469 = n1468 ^ x463;
  assign n1470 = n1469 ^ x464;
  assign n1471 = ~n1125 & n1470;
  assign n1472 = n1471 ^ x464;
  assign n1473 = n1472 ^ x465;
  assign n1474 = ~n1124 & ~n1473;
  assign n1475 = n1474 ^ x337;
  assign n1476 = n1475 ^ x466;
  assign n1477 = ~n1123 & n1476;
  assign n1478 = n1477 ^ x338;
  assign n1479 = n1478 ^ x467;
  assign n1480 = ~n1122 & ~n1479;
  assign n1481 = n1480 ^ x467;
  assign n1482 = n1481 ^ x468;
  assign n1483 = ~n1121 & n1482;
  assign n1484 = n1483 ^ x468;
  assign n1485 = n1484 ^ x469;
  assign n1486 = ~n1120 & n1485;
  assign n1487 = n1486 ^ x469;
  assign n1488 = n1487 ^ x470;
  assign n1489 = ~n1119 & ~n1488;
  assign n1490 = n1489 ^ x342;
  assign n1491 = n1490 ^ x471;
  assign n1492 = ~n1118 & n1491;
  assign n1493 = n1492 ^ x343;
  assign n1494 = n1493 ^ x472;
  assign n1495 = ~n1117 & n1494;
  assign n1496 = n1495 ^ x344;
  assign n1497 = n1496 ^ x473;
  assign n1498 = ~n1116 & n1497;
  assign n1499 = n1498 ^ x345;
  assign n1500 = n1499 ^ x474;
  assign n1501 = ~n1115 & ~n1500;
  assign n1502 = n1501 ^ x474;
  assign n1503 = n1502 ^ x475;
  assign n1504 = ~n1114 & ~n1503;
  assign n1505 = n1504 ^ x347;
  assign n1506 = n1505 ^ x476;
  assign n1507 = ~n1113 & n1506;
  assign n1508 = n1507 ^ x348;
  assign n1509 = n1508 ^ x477;
  assign n1510 = ~n1112 & ~n1509;
  assign n1511 = n1510 ^ x477;
  assign n1512 = n1511 ^ x478;
  assign n1513 = ~n1111 & n1512;
  assign n1514 = n1513 ^ x478;
  assign n1515 = n1514 ^ x479;
  assign n1516 = ~n1110 & n1515;
  assign n1517 = n1516 ^ x479;
  assign n1518 = n1517 ^ x480;
  assign n1519 = ~n1109 & n1518;
  assign n1520 = n1519 ^ x480;
  assign n1521 = n1520 ^ x481;
  assign n1522 = ~n1108 & ~n1521;
  assign n1523 = n1522 ^ x353;
  assign n1524 = n1523 ^ x482;
  assign n1525 = ~n1107 & n1524;
  assign n1526 = n1525 ^ x354;
  assign n1527 = n1526 ^ x483;
  assign n1528 = ~n1106 & ~n1527;
  assign n1529 = n1528 ^ x483;
  assign n1530 = n1529 ^ x484;
  assign n1531 = ~n1105 & n1530;
  assign n1532 = n1531 ^ x484;
  assign n1533 = n1532 ^ x485;
  assign n1534 = ~n1104 & n1533;
  assign n1535 = n1534 ^ x485;
  assign n1536 = n1535 ^ x486;
  assign n1537 = ~n1103 & ~n1536;
  assign n1538 = n1537 ^ x358;
  assign n1539 = n1538 ^ x487;
  assign n1540 = ~n1102 & n1539;
  assign n1541 = n1540 ^ x359;
  assign n1542 = n1541 ^ x488;
  assign n1543 = ~n1101 & n1542;
  assign n1544 = n1543 ^ x360;
  assign n1545 = n1544 ^ x489;
  assign n1546 = ~n1100 & n1545;
  assign n1547 = n1546 ^ x361;
  assign n1548 = n1547 ^ x490;
  assign n1549 = ~n1099 & n1548;
  assign n1550 = n1549 ^ x362;
  assign n1551 = n1550 ^ x491;
  assign n1552 = ~n1098 & n1551;
  assign n1553 = n1552 ^ x363;
  assign n1554 = n1553 ^ x492;
  assign n1555 = ~n1097 & ~n1554;
  assign n1556 = n1555 ^ x492;
  assign n1557 = n1556 ^ x493;
  assign n1558 = ~n1096 & ~n1557;
  assign n1559 = n1558 ^ x365;
  assign n1560 = n1559 ^ x494;
  assign n1561 = ~n1095 & n1560;
  assign n1562 = n1561 ^ x366;
  assign n1563 = n1562 ^ x495;
  assign n1564 = ~n1094 & ~n1563;
  assign n1565 = n1564 ^ x495;
  assign n1566 = n1565 ^ x496;
  assign n1567 = ~n1093 & n1566;
  assign n1568 = n1567 ^ x496;
  assign n1569 = n1568 ^ x497;
  assign n1570 = ~n1092 & n1569;
  assign n1571 = n1570 ^ x497;
  assign n1572 = n1571 ^ x498;
  assign n1573 = ~n1091 & n1572;
  assign n1574 = n1573 ^ x498;
  assign n1575 = n1574 ^ x499;
  assign n1576 = ~n1090 & ~n1575;
  assign n1577 = n1576 ^ x371;
  assign n1578 = n1577 ^ x500;
  assign n1579 = ~n1089 & n1578;
  assign n1580 = n1579 ^ x372;
  assign n1581 = n1580 ^ x501;
  assign n1582 = ~n1088 & ~n1581;
  assign n1583 = n1582 ^ x501;
  assign n1584 = n1583 ^ x502;
  assign n1585 = ~n1087 & ~n1584;
  assign n1586 = n1585 ^ x374;
  assign n1587 = n1586 ^ x503;
  assign n1588 = ~n1086 & n1587;
  assign n1589 = n1588 ^ x375;
  assign n1590 = n1589 ^ x504;
  assign n1591 = ~n1085 & ~n1590;
  assign n1592 = n1591 ^ x504;
  assign n1593 = n1592 ^ x505;
  assign n1594 = ~n1084 & n1593;
  assign n1595 = n1594 ^ x505;
  assign n1596 = n1595 ^ x506;
  assign n1597 = ~n1083 & n1596;
  assign n1598 = n1597 ^ x506;
  assign n1599 = ~n1082 & n1598;
  assign n1600 = n1081 & ~n1599;
  assign n1601 = n1600 ^ x511;
  assign n1602 = n1601 ^ x511;
  assign n1603 = n1074 & ~n1602;
  assign n1604 = n1603 ^ x511;
  assign n1605 = ~n1064 & n1604;
  assign n1606 = n1605 ^ x383;
  assign n1607 = n1063 & n1606;
  assign n1608 = n1607 ^ x382;
  assign n2660 = n1608 ^ n514;
  assign n516 = x254 ^ x126;
  assign n517 = x255 ^ x127;
  assign n518 = x253 ^ x125;
  assign n519 = x124 & ~x252;
  assign n520 = n519 ^ x253;
  assign n521 = ~n518 & ~n520;
  assign n522 = n521 ^ x253;
  assign n523 = n522 ^ x254;
  assign n524 = ~n516 & n523;
  assign n525 = n524 ^ x254;
  assign n526 = n525 ^ x255;
  assign n527 = n526 ^ x255;
  assign n528 = ~x125 & x253;
  assign n529 = ~x126 & x254;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~x123 & x251;
  assign n532 = ~x124 & x252;
  assign n533 = ~n531 & ~n532;
  assign n534 = n530 & n533;
  assign n535 = x123 & ~x251;
  assign n536 = x250 ^ x122;
  assign n537 = x249 ^ x121;
  assign n538 = x248 ^ x120;
  assign n539 = x247 ^ x119;
  assign n540 = x246 ^ x118;
  assign n541 = x245 ^ x117;
  assign n542 = x244 ^ x116;
  assign n543 = x243 ^ x115;
  assign n544 = x242 ^ x114;
  assign n545 = x241 ^ x113;
  assign n546 = x240 ^ x112;
  assign n547 = x239 ^ x111;
  assign n548 = x238 ^ x110;
  assign n549 = x237 ^ x109;
  assign n550 = x236 ^ x108;
  assign n551 = x235 ^ x107;
  assign n552 = x234 ^ x106;
  assign n553 = x233 ^ x105;
  assign n554 = x232 ^ x104;
  assign n555 = x231 ^ x103;
  assign n556 = x230 ^ x102;
  assign n557 = x229 ^ x101;
  assign n558 = x228 ^ x100;
  assign n559 = x227 ^ x99;
  assign n560 = x226 ^ x98;
  assign n561 = x225 ^ x97;
  assign n562 = x224 ^ x96;
  assign n563 = x223 ^ x95;
  assign n564 = x222 ^ x94;
  assign n565 = x221 ^ x93;
  assign n566 = x220 ^ x92;
  assign n567 = x219 ^ x91;
  assign n568 = x218 ^ x90;
  assign n569 = x217 ^ x89;
  assign n570 = x216 ^ x88;
  assign n571 = x215 ^ x87;
  assign n572 = x214 ^ x86;
  assign n573 = x213 ^ x85;
  assign n574 = x212 ^ x84;
  assign n575 = x211 ^ x83;
  assign n576 = x210 ^ x82;
  assign n577 = x209 ^ x81;
  assign n578 = x80 & ~x208;
  assign n579 = n578 ^ x209;
  assign n580 = n579 ^ x209;
  assign n581 = ~x70 & x198;
  assign n582 = ~x69 & x197;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~x68 & x196;
  assign n585 = n583 & ~n584;
  assign n586 = x195 ^ x67;
  assign n587 = x194 ^ x66;
  assign n588 = x193 ^ x65;
  assign n589 = x192 ^ x64;
  assign n590 = ~x63 & x191;
  assign n591 = n590 ^ x192;
  assign n592 = n591 ^ x192;
  assign n593 = ~x62 & x190;
  assign n594 = ~x61 & x189;
  assign n595 = ~n593 & ~n594;
  assign n596 = ~x59 & x187;
  assign n597 = ~x60 & x188;
  assign n598 = ~n596 & ~n597;
  assign n599 = n595 & n598;
  assign n600 = x59 & ~x187;
  assign n601 = x186 ^ x58;
  assign n602 = x185 ^ x57;
  assign n603 = x184 ^ x56;
  assign n604 = x183 ^ x55;
  assign n605 = x182 ^ x54;
  assign n606 = x181 ^ x53;
  assign n607 = x180 ^ x52;
  assign n608 = x179 ^ x51;
  assign n609 = x178 ^ x50;
  assign n610 = x177 ^ x49;
  assign n611 = x48 & ~x176;
  assign n612 = n611 ^ x177;
  assign n613 = n612 ^ x177;
  assign n614 = x39 & ~x167;
  assign n615 = x166 ^ x38;
  assign n616 = x165 ^ x37;
  assign n617 = x164 ^ x36;
  assign n618 = x163 ^ x35;
  assign n619 = x162 ^ x34;
  assign n620 = x161 ^ x33;
  assign n621 = x160 ^ x32;
  assign n622 = x159 ^ x31;
  assign n623 = x158 ^ x30;
  assign n624 = x157 ^ x29;
  assign n625 = x156 ^ x28;
  assign n626 = x155 ^ x27;
  assign n627 = x154 ^ x26;
  assign n628 = x153 ^ x25;
  assign n629 = x152 ^ x24;
  assign n630 = x151 ^ x23;
  assign n631 = x150 ^ x22;
  assign n632 = x149 ^ x21;
  assign n633 = x148 ^ x20;
  assign n634 = x147 ^ x19;
  assign n635 = x146 ^ x18;
  assign n636 = x145 ^ x17;
  assign n637 = x144 ^ x16;
  assign n638 = x143 ^ x15;
  assign n639 = x142 ^ x14;
  assign n640 = x141 ^ x13;
  assign n641 = x140 ^ x12;
  assign n642 = x139 ^ x11;
  assign n643 = x138 ^ x10;
  assign n644 = x137 ^ x9;
  assign n645 = x136 ^ x8;
  assign n646 = x135 ^ x7;
  assign n647 = x134 ^ x6;
  assign n648 = x133 ^ x5;
  assign n649 = x132 ^ x4;
  assign n650 = x131 ^ x3;
  assign n651 = x130 ^ x2;
  assign n652 = x129 ^ x1;
  assign n653 = x0 & ~x128;
  assign n654 = n653 ^ x129;
  assign n655 = ~n652 & ~n654;
  assign n656 = n655 ^ x129;
  assign n657 = n656 ^ x130;
  assign n658 = ~n651 & n657;
  assign n659 = n658 ^ x130;
  assign n660 = n659 ^ x131;
  assign n661 = ~n650 & n660;
  assign n662 = n661 ^ x131;
  assign n663 = n662 ^ x132;
  assign n664 = ~n649 & ~n663;
  assign n665 = n664 ^ x4;
  assign n666 = n665 ^ x133;
  assign n667 = ~n648 & n666;
  assign n668 = n667 ^ x5;
  assign n669 = n668 ^ x134;
  assign n670 = ~n647 & ~n669;
  assign n671 = n670 ^ x134;
  assign n672 = n671 ^ x135;
  assign n673 = ~n646 & ~n672;
  assign n674 = n673 ^ x7;
  assign n675 = n674 ^ x136;
  assign n676 = ~n645 & n675;
  assign n677 = n676 ^ x8;
  assign n678 = n677 ^ x137;
  assign n679 = ~n644 & ~n678;
  assign n680 = n679 ^ x137;
  assign n681 = n680 ^ x138;
  assign n682 = ~n643 & ~n681;
  assign n683 = n682 ^ x10;
  assign n684 = n683 ^ x139;
  assign n685 = ~n642 & n684;
  assign n686 = n685 ^ x11;
  assign n687 = n686 ^ x140;
  assign n688 = ~n641 & n687;
  assign n689 = n688 ^ x12;
  assign n690 = n689 ^ x141;
  assign n691 = ~n640 & n690;
  assign n692 = n691 ^ x13;
  assign n693 = n692 ^ x142;
  assign n694 = ~n639 & n693;
  assign n695 = n694 ^ x14;
  assign n696 = n695 ^ x143;
  assign n697 = ~n638 & n696;
  assign n698 = n697 ^ x15;
  assign n699 = n698 ^ x144;
  assign n700 = ~n637 & ~n699;
  assign n701 = n700 ^ x144;
  assign n702 = n701 ^ x145;
  assign n703 = ~n636 & ~n702;
  assign n704 = n703 ^ x17;
  assign n705 = n704 ^ x146;
  assign n706 = ~n635 & n705;
  assign n707 = n706 ^ x18;
  assign n708 = n707 ^ x147;
  assign n709 = ~n634 & ~n708;
  assign n710 = n709 ^ x147;
  assign n711 = n710 ^ x148;
  assign n712 = ~n633 & n711;
  assign n713 = n712 ^ x148;
  assign n714 = n713 ^ x149;
  assign n715 = ~n632 & n714;
  assign n716 = n715 ^ x149;
  assign n717 = n716 ^ x150;
  assign n718 = ~n631 & n717;
  assign n719 = n718 ^ x150;
  assign n720 = n719 ^ x151;
  assign n721 = ~n630 & n720;
  assign n722 = n721 ^ x151;
  assign n723 = n722 ^ x152;
  assign n724 = ~n629 & n723;
  assign n725 = n724 ^ x152;
  assign n726 = n725 ^ x153;
  assign n727 = ~n628 & ~n726;
  assign n728 = n727 ^ x25;
  assign n729 = n728 ^ x154;
  assign n730 = ~n627 & n729;
  assign n731 = n730 ^ x26;
  assign n732 = n731 ^ x155;
  assign n733 = ~n626 & ~n732;
  assign n734 = n733 ^ x155;
  assign n735 = n734 ^ x156;
  assign n736 = ~n625 & ~n735;
  assign n737 = n736 ^ x28;
  assign n738 = n737 ^ x157;
  assign n739 = ~n624 & n738;
  assign n740 = n739 ^ x29;
  assign n741 = n740 ^ x158;
  assign n742 = ~n623 & ~n741;
  assign n743 = n742 ^ x158;
  assign n744 = n743 ^ x159;
  assign n745 = ~n622 & ~n744;
  assign n746 = n745 ^ x31;
  assign n747 = n746 ^ x160;
  assign n748 = ~n621 & n747;
  assign n749 = n748 ^ x32;
  assign n750 = n749 ^ x161;
  assign n751 = ~n620 & ~n750;
  assign n752 = n751 ^ x161;
  assign n753 = n752 ^ x162;
  assign n754 = ~n619 & n753;
  assign n755 = n754 ^ x162;
  assign n756 = n755 ^ x163;
  assign n757 = ~n618 & n756;
  assign n758 = n757 ^ x163;
  assign n759 = n758 ^ x164;
  assign n760 = ~n617 & n759;
  assign n761 = n760 ^ x164;
  assign n762 = n761 ^ x165;
  assign n763 = ~n616 & ~n762;
  assign n764 = n763 ^ x37;
  assign n765 = n764 ^ x166;
  assign n766 = ~n615 & n765;
  assign n767 = n766 ^ x38;
  assign n768 = ~n614 & ~n767;
  assign n769 = ~x41 & x169;
  assign n770 = ~x42 & x170;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~x39 & x167;
  assign n773 = ~x40 & x168;
  assign n774 = ~n772 & ~n773;
  assign n775 = n771 & n774;
  assign n776 = ~n768 & n775;
  assign n777 = x43 & ~x171;
  assign n778 = x170 ^ x42;
  assign n779 = x169 ^ x41;
  assign n780 = x40 & ~x168;
  assign n781 = n780 ^ x169;
  assign n782 = ~n779 & ~n781;
  assign n783 = n782 ^ x169;
  assign n784 = n783 ^ x170;
  assign n785 = ~n778 & n784;
  assign n786 = n785 ^ x170;
  assign n787 = ~n777 & n786;
  assign n788 = ~n776 & n787;
  assign n789 = ~x46 & x174;
  assign n790 = ~x45 & x173;
  assign n791 = ~n789 & ~n790;
  assign n792 = ~x43 & x171;
  assign n793 = ~x44 & x172;
  assign n794 = ~n792 & ~n793;
  assign n795 = n791 & n794;
  assign n796 = ~n788 & n795;
  assign n797 = x47 & ~x175;
  assign n798 = x174 ^ x46;
  assign n799 = x173 ^ x45;
  assign n800 = x44 & ~x172;
  assign n801 = n800 ^ x173;
  assign n802 = ~n799 & ~n801;
  assign n803 = n802 ^ x173;
  assign n804 = n803 ^ x174;
  assign n805 = ~n798 & n804;
  assign n806 = n805 ^ x174;
  assign n807 = ~n797 & n806;
  assign n808 = ~n796 & n807;
  assign n809 = ~x48 & x176;
  assign n810 = ~x47 & x175;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n808 & n811;
  assign n813 = n812 ^ x177;
  assign n814 = n813 ^ x177;
  assign n815 = ~n613 & ~n814;
  assign n816 = n815 ^ x177;
  assign n817 = ~n610 & ~n816;
  assign n818 = n817 ^ x49;
  assign n819 = n818 ^ x178;
  assign n820 = ~n609 & ~n819;
  assign n821 = n820 ^ x178;
  assign n822 = n821 ^ x179;
  assign n823 = ~n608 & n822;
  assign n824 = n823 ^ x179;
  assign n825 = n824 ^ x180;
  assign n826 = ~n607 & n825;
  assign n827 = n826 ^ x180;
  assign n828 = n827 ^ x181;
  assign n829 = ~n606 & n828;
  assign n830 = n829 ^ x181;
  assign n831 = n830 ^ x182;
  assign n832 = ~n605 & n831;
  assign n833 = n832 ^ x182;
  assign n834 = n833 ^ x183;
  assign n835 = ~n604 & ~n834;
  assign n836 = n835 ^ x55;
  assign n837 = n836 ^ x184;
  assign n838 = ~n603 & n837;
  assign n839 = n838 ^ x56;
  assign n840 = n839 ^ x185;
  assign n841 = ~n602 & ~n840;
  assign n842 = n841 ^ x185;
  assign n843 = n842 ^ x186;
  assign n844 = ~n601 & n843;
  assign n845 = n844 ^ x186;
  assign n846 = ~n600 & n845;
  assign n847 = n599 & ~n846;
  assign n848 = x63 & ~x191;
  assign n849 = x190 ^ x62;
  assign n850 = x189 ^ x61;
  assign n851 = x60 & ~x188;
  assign n852 = n851 ^ x189;
  assign n853 = ~n850 & ~n852;
  assign n854 = n853 ^ x189;
  assign n855 = n854 ^ x190;
  assign n856 = ~n849 & n855;
  assign n857 = n856 ^ x190;
  assign n858 = ~n848 & n857;
  assign n859 = ~n847 & n858;
  assign n860 = n859 ^ x192;
  assign n861 = n860 ^ x192;
  assign n862 = ~n592 & ~n861;
  assign n863 = n862 ^ x192;
  assign n864 = ~n589 & n863;
  assign n865 = n864 ^ x64;
  assign n866 = n865 ^ x193;
  assign n867 = ~n588 & ~n866;
  assign n868 = n867 ^ x193;
  assign n869 = n868 ^ x194;
  assign n870 = ~n587 & ~n869;
  assign n871 = n870 ^ x66;
  assign n872 = n871 ^ x195;
  assign n873 = ~n586 & n872;
  assign n874 = n873 ^ x67;
  assign n875 = n585 & n874;
  assign n876 = x71 & ~x199;
  assign n877 = x198 ^ x70;
  assign n878 = x197 ^ x69;
  assign n879 = x68 & ~x196;
  assign n880 = n879 ^ x197;
  assign n881 = ~n878 & ~n880;
  assign n882 = n881 ^ x197;
  assign n883 = n882 ^ x198;
  assign n884 = ~n877 & n883;
  assign n885 = n884 ^ x198;
  assign n886 = ~n876 & n885;
  assign n887 = ~n875 & n886;
  assign n888 = ~x72 & x200;
  assign n889 = ~x71 & x199;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~n887 & n890;
  assign n892 = x73 & ~x201;
  assign n893 = x72 & ~x200;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n891 & n894;
  assign n896 = ~x74 & x202;
  assign n897 = ~x73 & x201;
  assign n898 = ~n896 & ~n897;
  assign n899 = ~n895 & n898;
  assign n900 = x75 & ~x203;
  assign n901 = x74 & ~x202;
  assign n902 = ~n900 & ~n901;
  assign n903 = ~n899 & n902;
  assign n904 = ~x76 & x204;
  assign n905 = ~x75 & x203;
  assign n906 = ~n904 & ~n905;
  assign n907 = ~n903 & n906;
  assign n908 = x77 & ~x205;
  assign n909 = x76 & ~x204;
  assign n910 = ~n908 & ~n909;
  assign n911 = ~n907 & n910;
  assign n912 = ~x78 & x206;
  assign n913 = ~x77 & x205;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~n911 & n914;
  assign n916 = x79 & ~x207;
  assign n917 = x78 & ~x206;
  assign n918 = ~n916 & ~n917;
  assign n919 = ~n915 & n918;
  assign n920 = ~x80 & x208;
  assign n921 = ~x79 & x207;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n919 & n922;
  assign n924 = n923 ^ x209;
  assign n925 = n924 ^ x209;
  assign n926 = ~n580 & ~n925;
  assign n927 = n926 ^ x209;
  assign n928 = ~n577 & ~n927;
  assign n929 = n928 ^ x81;
  assign n930 = n929 ^ x210;
  assign n931 = ~n576 & ~n930;
  assign n932 = n931 ^ x210;
  assign n933 = n932 ^ x211;
  assign n934 = ~n575 & n933;
  assign n935 = n934 ^ x211;
  assign n936 = n935 ^ x212;
  assign n937 = ~n574 & n936;
  assign n938 = n937 ^ x212;
  assign n939 = n938 ^ x213;
  assign n940 = ~n573 & n939;
  assign n941 = n940 ^ x213;
  assign n942 = n941 ^ x214;
  assign n943 = ~n572 & n942;
  assign n944 = n943 ^ x214;
  assign n945 = n944 ^ x215;
  assign n946 = ~n571 & n945;
  assign n947 = n946 ^ x215;
  assign n948 = n947 ^ x216;
  assign n949 = ~n570 & n948;
  assign n950 = n949 ^ x216;
  assign n951 = n950 ^ x217;
  assign n952 = ~n569 & ~n951;
  assign n953 = n952 ^ x89;
  assign n954 = n953 ^ x218;
  assign n955 = ~n568 & n954;
  assign n956 = n955 ^ x90;
  assign n957 = n956 ^ x219;
  assign n958 = ~n567 & n957;
  assign n959 = n958 ^ x91;
  assign n960 = n959 ^ x220;
  assign n961 = ~n566 & n960;
  assign n962 = n961 ^ x92;
  assign n963 = n962 ^ x221;
  assign n964 = ~n565 & n963;
  assign n965 = n964 ^ x93;
  assign n966 = n965 ^ x222;
  assign n967 = ~n564 & n966;
  assign n968 = n967 ^ x94;
  assign n969 = n968 ^ x223;
  assign n970 = ~n563 & ~n969;
  assign n971 = n970 ^ x223;
  assign n972 = n971 ^ x224;
  assign n973 = ~n562 & ~n972;
  assign n974 = n973 ^ x96;
  assign n975 = n974 ^ x225;
  assign n976 = ~n561 & n975;
  assign n977 = n976 ^ x97;
  assign n978 = n977 ^ x226;
  assign n979 = ~n560 & ~n978;
  assign n980 = n979 ^ x226;
  assign n981 = n980 ^ x227;
  assign n982 = ~n559 & n981;
  assign n983 = n982 ^ x227;
  assign n984 = n983 ^ x228;
  assign n985 = ~n558 & ~n984;
  assign n986 = n985 ^ x100;
  assign n987 = n986 ^ x229;
  assign n988 = ~n557 & n987;
  assign n989 = n988 ^ x101;
  assign n990 = n989 ^ x230;
  assign n991 = ~n556 & ~n990;
  assign n992 = n991 ^ x230;
  assign n993 = n992 ^ x231;
  assign n994 = ~n555 & n993;
  assign n995 = n994 ^ x231;
  assign n996 = n995 ^ x232;
  assign n997 = ~n554 & ~n996;
  assign n998 = n997 ^ x104;
  assign n999 = n998 ^ x233;
  assign n1000 = ~n553 & n999;
  assign n1001 = n1000 ^ x105;
  assign n1002 = n1001 ^ x234;
  assign n1003 = ~n552 & ~n1002;
  assign n1004 = n1003 ^ x234;
  assign n1005 = n1004 ^ x235;
  assign n1006 = ~n551 & n1005;
  assign n1007 = n1006 ^ x235;
  assign n1008 = n1007 ^ x236;
  assign n1009 = ~n550 & ~n1008;
  assign n1010 = n1009 ^ x108;
  assign n1011 = n1010 ^ x237;
  assign n1012 = ~n549 & n1011;
  assign n1013 = n1012 ^ x109;
  assign n1014 = n1013 ^ x238;
  assign n1015 = ~n548 & ~n1014;
  assign n1016 = n1015 ^ x238;
  assign n1017 = n1016 ^ x239;
  assign n1018 = ~n547 & n1017;
  assign n1019 = n1018 ^ x239;
  assign n1020 = n1019 ^ x240;
  assign n1021 = ~n546 & ~n1020;
  assign n1022 = n1021 ^ x112;
  assign n1023 = n1022 ^ x241;
  assign n1024 = ~n545 & n1023;
  assign n1025 = n1024 ^ x113;
  assign n1026 = n1025 ^ x242;
  assign n1027 = ~n544 & ~n1026;
  assign n1028 = n1027 ^ x242;
  assign n1029 = n1028 ^ x243;
  assign n1030 = ~n543 & ~n1029;
  assign n1031 = n1030 ^ x115;
  assign n1032 = n1031 ^ x244;
  assign n1033 = ~n542 & n1032;
  assign n1034 = n1033 ^ x116;
  assign n1035 = n1034 ^ x245;
  assign n1036 = ~n541 & ~n1035;
  assign n1037 = n1036 ^ x245;
  assign n1038 = n1037 ^ x246;
  assign n1039 = ~n540 & ~n1038;
  assign n1040 = n1039 ^ x118;
  assign n1041 = n1040 ^ x247;
  assign n1042 = ~n539 & n1041;
  assign n1043 = n1042 ^ x119;
  assign n1044 = n1043 ^ x248;
  assign n1045 = ~n538 & n1044;
  assign n1046 = n1045 ^ x120;
  assign n1047 = n1046 ^ x249;
  assign n1048 = ~n537 & n1047;
  assign n1049 = n1048 ^ x121;
  assign n1050 = n1049 ^ x250;
  assign n1051 = ~n536 & ~n1050;
  assign n1052 = n1051 ^ x250;
  assign n1053 = ~n535 & n1052;
  assign n1054 = n534 & ~n1053;
  assign n1055 = n1054 ^ x255;
  assign n1056 = n1055 ^ x255;
  assign n1057 = n527 & ~n1056;
  assign n1058 = n1057 ^ x255;
  assign n1059 = ~n517 & n1058;
  assign n1060 = n1059 ^ x127;
  assign n1061 = n516 & n1060;
  assign n1062 = n1061 ^ x126;
  assign n1609 = n1608 ^ n1062;
  assign n1612 = n518 & n1060;
  assign n1613 = n1612 ^ x125;
  assign n1610 = n1065 & n1606;
  assign n1611 = n1610 ^ x381;
  assign n1614 = n1613 ^ n1611;
  assign n1618 = x252 ^ x124;
  assign n1619 = n1060 & n1618;
  assign n1620 = n1619 ^ x124;
  assign n1615 = x508 ^ x380;
  assign n1616 = n1606 & n1615;
  assign n1617 = n1616 ^ x380;
  assign n1621 = n1620 ^ n1617;
  assign n1625 = x251 ^ x123;
  assign n1626 = n1060 & n1625;
  assign n1627 = n1626 ^ x123;
  assign n1622 = x507 ^ x379;
  assign n1623 = n1606 & n1622;
  assign n1624 = n1623 ^ x379;
  assign n1628 = n1627 ^ n1624;
  assign n1631 = n536 & n1060;
  assign n1632 = n1631 ^ x122;
  assign n1629 = n1083 & n1606;
  assign n1630 = n1629 ^ x378;
  assign n1633 = n1632 ^ n1630;
  assign n1636 = n537 & n1060;
  assign n1637 = n1636 ^ x121;
  assign n1634 = n1084 & n1606;
  assign n1635 = n1634 ^ x377;
  assign n1638 = n1637 ^ n1635;
  assign n1641 = n1085 & n1606;
  assign n1642 = n1641 ^ x376;
  assign n1639 = n538 & n1060;
  assign n1640 = n1639 ^ x120;
  assign n1643 = n1642 ^ n1640;
  assign n1646 = n539 & n1060;
  assign n1647 = n1646 ^ x119;
  assign n1644 = n1086 & n1606;
  assign n1645 = n1644 ^ x375;
  assign n1648 = n1647 ^ n1645;
  assign n1651 = n540 & n1060;
  assign n1652 = n1651 ^ x118;
  assign n1649 = n1087 & n1606;
  assign n1650 = n1649 ^ x374;
  assign n1653 = n1652 ^ n1650;
  assign n1656 = n541 & n1060;
  assign n1657 = n1656 ^ x117;
  assign n1654 = n1088 & n1606;
  assign n1655 = n1654 ^ x373;
  assign n1658 = n1657 ^ n1655;
  assign n1661 = n1089 & n1606;
  assign n1662 = n1661 ^ x372;
  assign n1659 = n542 & n1060;
  assign n1660 = n1659 ^ x116;
  assign n1663 = n1662 ^ n1660;
  assign n1666 = n1090 & n1606;
  assign n1667 = n1666 ^ x371;
  assign n1664 = n543 & n1060;
  assign n1665 = n1664 ^ x115;
  assign n1668 = n1667 ^ n1665;
  assign n1671 = n544 & n1060;
  assign n1672 = n1671 ^ x114;
  assign n1669 = n1091 & n1606;
  assign n1670 = n1669 ^ x370;
  assign n1673 = n1672 ^ n1670;
  assign n1676 = n545 & n1060;
  assign n1677 = n1676 ^ x113;
  assign n1674 = n1092 & n1606;
  assign n1675 = n1674 ^ x369;
  assign n1678 = n1677 ^ n1675;
  assign n1681 = n546 & n1060;
  assign n1682 = n1681 ^ x112;
  assign n1679 = n1093 & n1606;
  assign n1680 = n1679 ^ x368;
  assign n1683 = n1682 ^ n1680;
  assign n1686 = n547 & n1060;
  assign n1687 = n1686 ^ x111;
  assign n1684 = n1094 & n1606;
  assign n1685 = n1684 ^ x367;
  assign n1688 = n1687 ^ n1685;
  assign n1691 = n1095 & n1606;
  assign n1692 = n1691 ^ x366;
  assign n1689 = n548 & n1060;
  assign n1690 = n1689 ^ x110;
  assign n1693 = n1692 ^ n1690;
  assign n1696 = n1096 & n1606;
  assign n1697 = n1696 ^ x365;
  assign n1694 = n549 & n1060;
  assign n1695 = n1694 ^ x109;
  assign n1698 = n1697 ^ n1695;
  assign n1701 = n1097 & n1606;
  assign n1702 = n1701 ^ x364;
  assign n1699 = n550 & n1060;
  assign n1700 = n1699 ^ x108;
  assign n1703 = n1702 ^ n1700;
  assign n1706 = n551 & n1060;
  assign n1707 = n1706 ^ x107;
  assign n1704 = n1098 & n1606;
  assign n1705 = n1704 ^ x363;
  assign n1708 = n1707 ^ n1705;
  assign n1711 = n552 & n1060;
  assign n1712 = n1711 ^ x106;
  assign n1709 = n1099 & n1606;
  assign n1710 = n1709 ^ x362;
  assign n1713 = n1712 ^ n1710;
  assign n1716 = n553 & n1060;
  assign n1717 = n1716 ^ x105;
  assign n1714 = n1100 & n1606;
  assign n1715 = n1714 ^ x361;
  assign n1718 = n1717 ^ n1715;
  assign n1721 = n1101 & n1606;
  assign n1722 = n1721 ^ x360;
  assign n1719 = n554 & n1060;
  assign n1720 = n1719 ^ x104;
  assign n1723 = n1722 ^ n1720;
  assign n1726 = n1102 & n1606;
  assign n1727 = n1726 ^ x359;
  assign n1724 = n555 & n1060;
  assign n1725 = n1724 ^ x103;
  assign n1728 = n1727 ^ n1725;
  assign n1731 = n556 & n1060;
  assign n1732 = n1731 ^ x102;
  assign n1729 = n1103 & n1606;
  assign n1730 = n1729 ^ x358;
  assign n1733 = n1732 ^ n1730;
  assign n1736 = n1104 & n1606;
  assign n1737 = n1736 ^ x357;
  assign n1734 = n557 & n1060;
  assign n1735 = n1734 ^ x101;
  assign n1738 = n1737 ^ n1735;
  assign n1741 = n1105 & n1606;
  assign n1742 = n1741 ^ x356;
  assign n1739 = n558 & n1060;
  assign n1740 = n1739 ^ x100;
  assign n1743 = n1742 ^ n1740;
  assign n1746 = n559 & n1060;
  assign n1747 = n1746 ^ x99;
  assign n1744 = n1106 & n1606;
  assign n1745 = n1744 ^ x355;
  assign n1748 = n1747 ^ n1745;
  assign n1751 = n560 & n1060;
  assign n1752 = n1751 ^ x98;
  assign n1749 = n1107 & n1606;
  assign n1750 = n1749 ^ x354;
  assign n1753 = n1752 ^ n1750;
  assign n1756 = n1108 & n1606;
  assign n1757 = n1756 ^ x353;
  assign n1754 = n561 & n1060;
  assign n1755 = n1754 ^ x97;
  assign n1758 = n1757 ^ n1755;
  assign n1761 = n562 & n1060;
  assign n1762 = n1761 ^ x96;
  assign n1759 = n1109 & n1606;
  assign n1760 = n1759 ^ x352;
  assign n1763 = n1762 ^ n1760;
  assign n1766 = n563 & n1060;
  assign n1767 = n1766 ^ x95;
  assign n1764 = n1110 & n1606;
  assign n1765 = n1764 ^ x351;
  assign n1768 = n1767 ^ n1765;
  assign n1771 = n564 & n1060;
  assign n1772 = n1771 ^ x94;
  assign n1769 = n1111 & n1606;
  assign n1770 = n1769 ^ x350;
  assign n1773 = n1772 ^ n1770;
  assign n1776 = n565 & n1060;
  assign n1777 = n1776 ^ x93;
  assign n1774 = n1112 & n1606;
  assign n1775 = n1774 ^ x349;
  assign n1778 = n1777 ^ n1775;
  assign n1781 = n1113 & n1606;
  assign n1782 = n1781 ^ x348;
  assign n1779 = n566 & n1060;
  assign n1780 = n1779 ^ x92;
  assign n1783 = n1782 ^ n1780;
  assign n1786 = n1114 & n1606;
  assign n1787 = n1786 ^ x347;
  assign n1784 = n567 & n1060;
  assign n1785 = n1784 ^ x91;
  assign n1788 = n1787 ^ n1785;
  assign n1791 = n1115 & n1606;
  assign n1792 = n1791 ^ x346;
  assign n1789 = n568 & n1060;
  assign n1790 = n1789 ^ x90;
  assign n1793 = n1792 ^ n1790;
  assign n1796 = n569 & n1060;
  assign n1797 = n1796 ^ x89;
  assign n1794 = n1116 & n1606;
  assign n1795 = n1794 ^ x345;
  assign n1798 = n1797 ^ n1795;
  assign n1801 = n1117 & n1606;
  assign n1802 = n1801 ^ x344;
  assign n1799 = n570 & n1060;
  assign n1800 = n1799 ^ x88;
  assign n1803 = n1802 ^ n1800;
  assign n1806 = n1118 & n1606;
  assign n1807 = n1806 ^ x343;
  assign n1804 = n571 & n1060;
  assign n1805 = n1804 ^ x87;
  assign n1808 = n1807 ^ n1805;
  assign n1811 = n1119 & n1606;
  assign n1812 = n1811 ^ x342;
  assign n1809 = n572 & n1060;
  assign n1810 = n1809 ^ x86;
  assign n1813 = n1812 ^ n1810;
  assign n1816 = n1120 & n1606;
  assign n1817 = n1816 ^ x341;
  assign n1814 = n573 & n1060;
  assign n1815 = n1814 ^ x85;
  assign n1818 = n1817 ^ n1815;
  assign n1821 = n574 & n1060;
  assign n1822 = n1821 ^ x84;
  assign n1819 = n1121 & n1606;
  assign n1820 = n1819 ^ x340;
  assign n1823 = n1822 ^ n1820;
  assign n1826 = n1122 & n1606;
  assign n1827 = n1826 ^ x339;
  assign n1824 = n575 & n1060;
  assign n1825 = n1824 ^ x83;
  assign n1828 = n1827 ^ n1825;
  assign n1831 = n576 & n1060;
  assign n1832 = n1831 ^ x82;
  assign n1829 = n1123 & n1606;
  assign n1830 = n1829 ^ x338;
  assign n1833 = n1832 ^ n1830;
  assign n1836 = n1124 & n1606;
  assign n1837 = n1836 ^ x337;
  assign n1834 = n577 & n1060;
  assign n1835 = n1834 ^ x81;
  assign n1838 = n1837 ^ n1835;
  assign n1842 = n1125 & n1606;
  assign n1843 = n1842 ^ x336;
  assign n1839 = x208 ^ x80;
  assign n1840 = n1060 & n1839;
  assign n1841 = n1840 ^ x80;
  assign n1844 = n1843 ^ n1841;
  assign n1848 = n1126 & n1606;
  assign n1849 = n1848 ^ x335;
  assign n1845 = x207 ^ x79;
  assign n1846 = n1060 & n1845;
  assign n1847 = n1846 ^ x79;
  assign n1850 = n1849 ^ n1847;
  assign n1853 = x206 ^ x78;
  assign n1854 = n1060 & n1853;
  assign n1855 = n1854 ^ x78;
  assign n1851 = n1127 & n1606;
  assign n1852 = n1851 ^ x334;
  assign n1856 = n1855 ^ n1852;
  assign n1860 = n1128 & n1606;
  assign n1861 = n1860 ^ x333;
  assign n1857 = x205 ^ x77;
  assign n1858 = n1060 & n1857;
  assign n1859 = n1858 ^ x77;
  assign n1862 = n1861 ^ n1859;
  assign n1865 = x204 ^ x76;
  assign n1866 = n1060 & n1865;
  assign n1867 = n1866 ^ x76;
  assign n1863 = n1129 & n1606;
  assign n1864 = n1863 ^ x332;
  assign n1868 = n1867 ^ n1864;
  assign n1871 = x203 ^ x75;
  assign n1872 = n1060 & n1871;
  assign n1873 = n1872 ^ x75;
  assign n1869 = n1130 & n1606;
  assign n1870 = n1869 ^ x331;
  assign n1874 = n1873 ^ n1870;
  assign n1877 = x202 ^ x74;
  assign n1878 = n1060 & n1877;
  assign n1879 = n1878 ^ x74;
  assign n1875 = n1131 & n1606;
  assign n1876 = n1875 ^ x330;
  assign n1880 = n1879 ^ n1876;
  assign n1883 = x201 ^ x73;
  assign n1884 = n1060 & n1883;
  assign n1885 = n1884 ^ x73;
  assign n1881 = n1132 & n1606;
  assign n1882 = n1881 ^ x329;
  assign n1886 = n1885 ^ n1882;
  assign n1890 = n1133 & n1606;
  assign n1891 = n1890 ^ x328;
  assign n1887 = x200 ^ x72;
  assign n1888 = n1060 & n1887;
  assign n1889 = n1888 ^ x72;
  assign n1892 = n1891 ^ n1889;
  assign n1896 = x455 ^ x327;
  assign n1897 = n1606 & n1896;
  assign n1898 = n1897 ^ x327;
  assign n1893 = x199 ^ x71;
  assign n1894 = n1060 & n1893;
  assign n1895 = n1894 ^ x71;
  assign n1899 = n1898 ^ n1895;
  assign n1902 = n877 & n1060;
  assign n1903 = n1902 ^ x70;
  assign n1900 = n1432 & n1606;
  assign n1901 = n1900 ^ x326;
  assign n1904 = n1903 ^ n1901;
  assign n1907 = n1433 & n1606;
  assign n1908 = n1907 ^ x325;
  assign n1905 = n878 & n1060;
  assign n1906 = n1905 ^ x69;
  assign n1909 = n1908 ^ n1906;
  assign n1913 = x196 ^ x68;
  assign n1914 = n1060 & n1913;
  assign n1915 = n1914 ^ x68;
  assign n1910 = x452 ^ x324;
  assign n1911 = n1606 & n1910;
  assign n1912 = n1911 ^ x324;
  assign n1916 = n1915 ^ n1912;
  assign n1919 = x451 ^ x323;
  assign n1920 = n1606 & n1919;
  assign n1921 = n1920 ^ x323;
  assign n1917 = n586 & n1060;
  assign n1918 = n1917 ^ x67;
  assign n1922 = n1921 ^ n1918;
  assign n1925 = n1145 & n1606;
  assign n1926 = n1925 ^ x322;
  assign n1923 = n587 & n1060;
  assign n1924 = n1923 ^ x66;
  assign n1927 = n1926 ^ n1924;
  assign n1930 = n588 & n1060;
  assign n1931 = n1930 ^ x65;
  assign n1928 = n1146 & n1606;
  assign n1929 = n1928 ^ x321;
  assign n1932 = n1931 ^ n1929;
  assign n1935 = x448 ^ x320;
  assign n1936 = n1606 & n1935;
  assign n1937 = n1936 ^ x320;
  assign n1933 = n589 & n1060;
  assign n1934 = n1933 ^ x64;
  assign n1938 = n1937 ^ n1934;
  assign n1941 = x191 ^ x63;
  assign n1942 = n1060 & n1941;
  assign n1943 = n1942 ^ x63;
  assign n1939 = n1412 & n1606;
  assign n1940 = n1939 ^ x319;
  assign n1944 = n1943 ^ n1940;
  assign n1947 = x446 ^ x318;
  assign n1948 = n1606 & n1947;
  assign n1949 = n1948 ^ x318;
  assign n1945 = n849 & n1060;
  assign n1946 = n1945 ^ x62;
  assign n1950 = n1949 ^ n1946;
  assign n1953 = x445 ^ x317;
  assign n1954 = n1606 & n1953;
  assign n1955 = n1954 ^ x317;
  assign n1951 = n850 & n1060;
  assign n1952 = n1951 ^ x61;
  assign n1956 = n1955 ^ n1952;
  assign n1960 = x444 ^ x316;
  assign n1961 = n1606 & n1960;
  assign n1962 = n1961 ^ x316;
  assign n1957 = x188 ^ x60;
  assign n1958 = n1060 & n1957;
  assign n1959 = n1958 ^ x60;
  assign n1963 = n1962 ^ n1959;
  assign n1967 = x443 ^ x315;
  assign n1968 = n1606 & n1967;
  assign n1969 = n1968 ^ x315;
  assign n1964 = x187 ^ x59;
  assign n1965 = n1060 & n1964;
  assign n1966 = n1965 ^ x59;
  assign n1970 = n1969 ^ n1966;
  assign n1973 = n601 & n1060;
  assign n1974 = n1973 ^ x58;
  assign n1971 = n1151 & n1606;
  assign n1972 = n1971 ^ x314;
  assign n1975 = n1974 ^ n1972;
  assign n1978 = n602 & n1060;
  assign n1979 = n1978 ^ x57;
  assign n1976 = n1152 & n1606;
  assign n1977 = n1976 ^ x313;
  assign n1980 = n1979 ^ n1977;
  assign n1983 = n1153 & n1606;
  assign n1984 = n1983 ^ x312;
  assign n1981 = n603 & n1060;
  assign n1982 = n1981 ^ x56;
  assign n1985 = n1984 ^ n1982;
  assign n1988 = n1154 & n1606;
  assign n1989 = n1988 ^ x311;
  assign n1986 = n604 & n1060;
  assign n1987 = n1986 ^ x55;
  assign n1990 = n1989 ^ n1987;
  assign n1993 = n1155 & n1606;
  assign n1994 = n1993 ^ x310;
  assign n1991 = n605 & n1060;
  assign n1992 = n1991 ^ x54;
  assign n1995 = n1994 ^ n1992;
  assign n1998 = n606 & n1060;
  assign n1999 = n1998 ^ x53;
  assign n1996 = n1156 & n1606;
  assign n1997 = n1996 ^ x309;
  assign n2000 = n1999 ^ n1997;
  assign n2003 = n1157 & n1606;
  assign n2004 = n2003 ^ x308;
  assign n2001 = n607 & n1060;
  assign n2002 = n2001 ^ x52;
  assign n2005 = n2004 ^ n2002;
  assign n2009 = n608 & n1060;
  assign n2010 = n2009 ^ x51;
  assign n2006 = x435 ^ x307;
  assign n2007 = n1606 & n2006;
  assign n2008 = n2007 ^ x307;
  assign n2011 = n2010 ^ n2008;
  assign n2014 = x434 ^ x306;
  assign n2015 = n1606 & n2014;
  assign n2016 = n2015 ^ x306;
  assign n2012 = n609 & n1060;
  assign n2013 = n2012 ^ x50;
  assign n2017 = n2016 ^ n2013;
  assign n2020 = x433 ^ x305;
  assign n2021 = n1606 & n2020;
  assign n2022 = n2021 ^ x305;
  assign n2018 = n610 & n1060;
  assign n2019 = n2018 ^ x49;
  assign n2023 = n2022 ^ n2019;
  assign n2027 = x176 ^ x48;
  assign n2028 = n1060 & n2027;
  assign n2029 = n2028 ^ x48;
  assign n2024 = x432 ^ x304;
  assign n2025 = n1606 & n2024;
  assign n2026 = n2025 ^ x304;
  assign n2030 = n2029 ^ n2026;
  assign n2034 = x431 ^ x303;
  assign n2035 = n1606 & n2034;
  assign n2036 = n2035 ^ x303;
  assign n2031 = x175 ^ x47;
  assign n2032 = n1060 & n2031;
  assign n2033 = n2032 ^ x47;
  assign n2037 = n2036 ^ n2033;
  assign n2040 = n1345 & n1606;
  assign n2041 = n2040 ^ x302;
  assign n2038 = n798 & n1060;
  assign n2039 = n2038 ^ x46;
  assign n2042 = n2041 ^ n2039;
  assign n2045 = n1346 & n1606;
  assign n2046 = n2045 ^ x301;
  assign n2043 = n799 & n1060;
  assign n2044 = n2043 ^ x45;
  assign n2047 = n2046 ^ n2044;
  assign n2051 = x428 ^ x300;
  assign n2052 = n1606 & n2051;
  assign n2053 = n2052 ^ x300;
  assign n2048 = x172 ^ x44;
  assign n2049 = n1060 & n2048;
  assign n2050 = n2049 ^ x44;
  assign n2054 = n2053 ^ n2050;
  assign n2058 = x171 ^ x43;
  assign n2059 = n1060 & n2058;
  assign n2060 = n2059 ^ x43;
  assign n2055 = x427 ^ x299;
  assign n2056 = n1606 & n2055;
  assign n2057 = n2056 ^ x299;
  assign n2061 = n2060 ^ n2057;
  assign n2064 = n1325 & n1606;
  assign n2065 = n2064 ^ x298;
  assign n2062 = n778 & n1060;
  assign n2063 = n2062 ^ x42;
  assign n2066 = n2065 ^ n2063;
  assign n2069 = n1326 & n1606;
  assign n2070 = n2069 ^ x297;
  assign n2067 = n779 & n1060;
  assign n2068 = n2067 ^ x41;
  assign n2071 = n2070 ^ n2068;
  assign n2075 = x424 ^ x296;
  assign n2076 = n1606 & n2075;
  assign n2077 = n2076 ^ x296;
  assign n2072 = x168 ^ x40;
  assign n2073 = n1060 & n2072;
  assign n2074 = n2073 ^ x40;
  assign n2078 = n2077 ^ n2074;
  assign n2082 = x423 ^ x295;
  assign n2083 = n1606 & n2082;
  assign n2084 = n2083 ^ x295;
  assign n2079 = x167 ^ x39;
  assign n2080 = n1060 & n2079;
  assign n2081 = n2080 ^ x39;
  assign n2085 = n2084 ^ n2081;
  assign n2088 = n1169 & n1606;
  assign n2089 = n2088 ^ x294;
  assign n2086 = n615 & n1060;
  assign n2087 = n2086 ^ x38;
  assign n2090 = n2089 ^ n2087;
  assign n2093 = n616 & n1060;
  assign n2094 = n2093 ^ x37;
  assign n2091 = n1170 & n1606;
  assign n2092 = n2091 ^ x293;
  assign n2095 = n2094 ^ n2092;
  assign n2098 = n1171 & n1606;
  assign n2099 = n2098 ^ x292;
  assign n2096 = n617 & n1060;
  assign n2097 = n2096 ^ x36;
  assign n2100 = n2099 ^ n2097;
  assign n2103 = n618 & n1060;
  assign n2104 = n2103 ^ x35;
  assign n2101 = n1172 & n1606;
  assign n2102 = n2101 ^ x291;
  assign n2105 = n2104 ^ n2102;
  assign n2108 = n619 & n1060;
  assign n2109 = n2108 ^ x34;
  assign n2106 = n1173 & n1606;
  assign n2107 = n2106 ^ x290;
  assign n2110 = n2109 ^ n2107;
  assign n2113 = n1174 & n1606;
  assign n2114 = n2113 ^ x289;
  assign n2111 = n620 & n1060;
  assign n2112 = n2111 ^ x33;
  assign n2115 = n2114 ^ n2112;
  assign n2118 = n1175 & n1606;
  assign n2119 = n2118 ^ x288;
  assign n2116 = n621 & n1060;
  assign n2117 = n2116 ^ x32;
  assign n2120 = n2119 ^ n2117;
  assign n2123 = n1176 & n1606;
  assign n2124 = n2123 ^ x287;
  assign n2121 = n622 & n1060;
  assign n2122 = n2121 ^ x31;
  assign n2125 = n2124 ^ n2122;
  assign n2128 = n623 & n1060;
  assign n2129 = n2128 ^ x30;
  assign n2126 = n1177 & n1606;
  assign n2127 = n2126 ^ x286;
  assign n2130 = n2129 ^ n2127;
  assign n2133 = n1178 & n1606;
  assign n2134 = n2133 ^ x285;
  assign n2131 = n624 & n1060;
  assign n2132 = n2131 ^ x29;
  assign n2135 = n2134 ^ n2132;
  assign n2138 = n1179 & n1606;
  assign n2139 = n2138 ^ x284;
  assign n2136 = n625 & n1060;
  assign n2137 = n2136 ^ x28;
  assign n2140 = n2139 ^ n2137;
  assign n2143 = n626 & n1060;
  assign n2144 = n2143 ^ x27;
  assign n2141 = n1180 & n1606;
  assign n2142 = n2141 ^ x283;
  assign n2145 = n2144 ^ n2142;
  assign n2148 = n1181 & n1606;
  assign n2149 = n2148 ^ x282;
  assign n2146 = n627 & n1060;
  assign n2147 = n2146 ^ x26;
  assign n2150 = n2149 ^ n2147;
  assign n2153 = n1182 & n1606;
  assign n2154 = n2153 ^ x281;
  assign n2151 = n628 & n1060;
  assign n2152 = n2151 ^ x25;
  assign n2155 = n2154 ^ n2152;
  assign n2158 = n1183 & n1606;
  assign n2159 = n2158 ^ x280;
  assign n2156 = n629 & n1060;
  assign n2157 = n2156 ^ x24;
  assign n2160 = n2159 ^ n2157;
  assign n2163 = n1184 & n1606;
  assign n2164 = n2163 ^ x279;
  assign n2161 = n630 & n1060;
  assign n2162 = n2161 ^ x23;
  assign n2165 = n2164 ^ n2162;
  assign n2168 = n631 & n1060;
  assign n2169 = n2168 ^ x22;
  assign n2166 = n1185 & n1606;
  assign n2167 = n2166 ^ x278;
  assign n2170 = n2169 ^ n2167;
  assign n2173 = n632 & n1060;
  assign n2174 = n2173 ^ x21;
  assign n2171 = n1186 & n1606;
  assign n2172 = n2171 ^ x277;
  assign n2175 = n2174 ^ n2172;
  assign n2178 = n1187 & n1606;
  assign n2179 = n2178 ^ x276;
  assign n2176 = n633 & n1060;
  assign n2177 = n2176 ^ x20;
  assign n2180 = n2179 ^ n2177;
  assign n2183 = n634 & n1060;
  assign n2184 = n2183 ^ x19;
  assign n2181 = n1188 & n1606;
  assign n2182 = n2181 ^ x275;
  assign n2185 = n2184 ^ n2182;
  assign n2188 = n1189 & n1606;
  assign n2189 = n2188 ^ x274;
  assign n2186 = n635 & n1060;
  assign n2187 = n2186 ^ x18;
  assign n2190 = n2189 ^ n2187;
  assign n2193 = n1190 & n1606;
  assign n2194 = n2193 ^ x273;
  assign n2191 = n636 & n1060;
  assign n2192 = n2191 ^ x17;
  assign n2195 = n2194 ^ n2192;
  assign n2198 = n637 & n1060;
  assign n2199 = n2198 ^ x16;
  assign n2196 = n1191 & n1606;
  assign n2197 = n2196 ^ x272;
  assign n2200 = n2199 ^ n2197;
  assign n2203 = n1192 & n1606;
  assign n2204 = n2203 ^ x271;
  assign n2201 = n638 & n1060;
  assign n2202 = n2201 ^ x15;
  assign n2205 = n2204 ^ n2202;
  assign n2208 = n1193 & n1606;
  assign n2209 = n2208 ^ x270;
  assign n2206 = n639 & n1060;
  assign n2207 = n2206 ^ x14;
  assign n2210 = n2209 ^ n2207;
  assign n2213 = n640 & n1060;
  assign n2214 = n2213 ^ x13;
  assign n2211 = n1194 & n1606;
  assign n2212 = n2211 ^ x269;
  assign n2215 = n2214 ^ n2212;
  assign n2218 = n641 & n1060;
  assign n2219 = n2218 ^ x12;
  assign n2216 = n1195 & n1606;
  assign n2217 = n2216 ^ x268;
  assign n2220 = n2219 ^ n2217;
  assign n2223 = n1196 & n1606;
  assign n2224 = n2223 ^ x267;
  assign n2221 = n642 & n1060;
  assign n2222 = n2221 ^ x11;
  assign n2225 = n2224 ^ n2222;
  assign n2228 = n643 & n1060;
  assign n2229 = n2228 ^ x10;
  assign n2226 = n1197 & n1606;
  assign n2227 = n2226 ^ x266;
  assign n2230 = n2229 ^ n2227;
  assign n2233 = n644 & n1060;
  assign n2234 = n2233 ^ x9;
  assign n2231 = n1198 & n1606;
  assign n2232 = n2231 ^ x265;
  assign n2235 = n2234 ^ n2232;
  assign n2238 = n645 & n1060;
  assign n2239 = n2238 ^ x8;
  assign n2236 = n1199 & n1606;
  assign n2237 = n2236 ^ x264;
  assign n2240 = n2239 ^ n2237;
  assign n2243 = n1200 & n1606;
  assign n2244 = n2243 ^ x263;
  assign n2241 = n646 & n1060;
  assign n2242 = n2241 ^ x7;
  assign n2245 = n2244 ^ n2242;
  assign n2248 = n647 & n1060;
  assign n2249 = n2248 ^ x6;
  assign n2246 = n1201 & n1606;
  assign n2247 = n2246 ^ x262;
  assign n2250 = n2249 ^ n2247;
  assign n2253 = n1202 & n1606;
  assign n2254 = n2253 ^ x261;
  assign n2251 = n648 & n1060;
  assign n2252 = n2251 ^ x5;
  assign n2255 = n2254 ^ n2252;
  assign n2258 = n1203 & n1606;
  assign n2259 = n2258 ^ x260;
  assign n2256 = n649 & n1060;
  assign n2257 = n2256 ^ x4;
  assign n2260 = n2259 ^ n2257;
  assign n2263 = n1204 & n1606;
  assign n2264 = n2263 ^ x259;
  assign n2261 = n650 & n1060;
  assign n2262 = n2261 ^ x3;
  assign n2265 = n2264 ^ n2262;
  assign n2268 = n651 & n1060;
  assign n2269 = n2268 ^ x2;
  assign n2266 = n1205 & n1606;
  assign n2267 = n2266 ^ x258;
  assign n2270 = n2269 ^ n2267;
  assign n2273 = n652 & n1060;
  assign n2274 = n2273 ^ x1;
  assign n2271 = n1206 & n1606;
  assign n2272 = n2271 ^ x257;
  assign n2275 = n2274 ^ n2272;
  assign n2276 = x384 ^ x256;
  assign n2277 = n1606 & n2276;
  assign n2278 = n2277 ^ x256;
  assign n2279 = x128 ^ x0;
  assign n2280 = n1060 & n2279;
  assign n2281 = n2280 ^ x0;
  assign n2282 = ~n2278 & n2281;
  assign n2283 = n2282 ^ n2274;
  assign n2284 = ~n2275 & n2283;
  assign n2285 = n2284 ^ n2274;
  assign n2286 = n2285 ^ n2269;
  assign n2287 = ~n2270 & n2286;
  assign n2288 = n2287 ^ n2269;
  assign n2289 = n2288 ^ n2262;
  assign n2290 = ~n2265 & ~n2289;
  assign n2291 = n2290 ^ n2264;
  assign n2292 = n2291 ^ n2259;
  assign n2293 = ~n2260 & ~n2292;
  assign n2294 = n2293 ^ n2257;
  assign n2295 = n2294 ^ n2254;
  assign n2296 = ~n2255 & ~n2295;
  assign n2297 = n2296 ^ n2254;
  assign n2298 = n2297 ^ n2249;
  assign n2299 = ~n2250 & n2298;
  assign n2300 = n2299 ^ n2247;
  assign n2301 = n2300 ^ n2244;
  assign n2302 = ~n2245 & ~n2301;
  assign n2303 = n2302 ^ n2242;
  assign n2304 = n2303 ^ n2239;
  assign n2305 = ~n2240 & n2304;
  assign n2306 = n2305 ^ n2239;
  assign n2307 = n2306 ^ n2234;
  assign n2308 = ~n2235 & n2307;
  assign n2309 = n2308 ^ n2234;
  assign n2310 = n2309 ^ n2227;
  assign n2311 = ~n2230 & ~n2310;
  assign n2312 = n2311 ^ n2227;
  assign n2313 = n2312 ^ n2224;
  assign n2314 = ~n2225 & n2313;
  assign n2315 = n2314 ^ n2224;
  assign n2316 = n2315 ^ n2217;
  assign n2317 = ~n2220 & n2316;
  assign n2318 = n2317 ^ n2217;
  assign n2319 = n2318 ^ n2214;
  assign n2320 = ~n2215 & ~n2319;
  assign n2321 = n2320 ^ n2214;
  assign n2322 = n2321 ^ n2207;
  assign n2323 = ~n2210 & ~n2322;
  assign n2324 = n2323 ^ n2209;
  assign n2325 = n2324 ^ n2204;
  assign n2326 = ~n2205 & ~n2325;
  assign n2327 = n2326 ^ n2202;
  assign n2328 = n2327 ^ n2199;
  assign n2329 = ~n2200 & n2328;
  assign n2330 = n2329 ^ n2199;
  assign n2331 = n2330 ^ n2194;
  assign n2332 = ~n2195 & n2331;
  assign n2333 = n2332 ^ n2192;
  assign n2334 = n2333 ^ n2189;
  assign n2335 = ~n2190 & ~n2334;
  assign n2336 = n2335 ^ n2189;
  assign n2337 = n2336 ^ n2184;
  assign n2338 = ~n2185 & n2337;
  assign n2339 = n2338 ^ n2182;
  assign n2340 = n2339 ^ n2179;
  assign n2341 = ~n2180 & ~n2340;
  assign n2342 = n2341 ^ n2177;
  assign n2343 = n2342 ^ n2174;
  assign n2344 = ~n2175 & n2343;
  assign n2345 = n2344 ^ n2174;
  assign n2346 = n2345 ^ n2169;
  assign n2347 = ~n2170 & n2346;
  assign n2348 = n2347 ^ n2169;
  assign n2349 = n2348 ^ n2162;
  assign n2350 = ~n2165 & ~n2349;
  assign n2351 = n2350 ^ n2164;
  assign n2352 = n2351 ^ n2159;
  assign n2353 = ~n2160 & ~n2352;
  assign n2354 = n2353 ^ n2157;
  assign n2355 = n2354 ^ n2154;
  assign n2356 = ~n2155 & ~n2355;
  assign n2357 = n2356 ^ n2154;
  assign n2358 = n2357 ^ n2149;
  assign n2359 = ~n2150 & ~n2358;
  assign n2360 = n2359 ^ n2147;
  assign n2361 = n2360 ^ n2144;
  assign n2362 = ~n2145 & n2361;
  assign n2363 = n2362 ^ n2144;
  assign n2364 = n2363 ^ n2139;
  assign n2365 = ~n2140 & n2364;
  assign n2366 = n2365 ^ n2137;
  assign n2367 = n2366 ^ n2134;
  assign n2368 = ~n2135 & n2367;
  assign n2369 = n2368 ^ n2132;
  assign n2370 = n2369 ^ n2129;
  assign n2371 = ~n2130 & n2370;
  assign n2372 = n2371 ^ n2129;
  assign n2373 = n2372 ^ n2124;
  assign n2374 = ~n2125 & n2373;
  assign n2375 = n2374 ^ n2122;
  assign n2376 = n2375 ^ n2119;
  assign n2377 = ~n2120 & ~n2376;
  assign n2378 = n2377 ^ n2119;
  assign n2379 = n2378 ^ n2114;
  assign n2380 = ~n2115 & ~n2379;
  assign n2381 = n2380 ^ n2112;
  assign n2382 = n2381 ^ n2109;
  assign n2383 = ~n2110 & n2382;
  assign n2384 = n2383 ^ n2109;
  assign n2385 = n2384 ^ n2102;
  assign n2386 = ~n2105 & n2385;
  assign n2387 = n2386 ^ n2104;
  assign n2388 = n2387 ^ n2099;
  assign n2389 = ~n2100 & n2388;
  assign n2390 = n2389 ^ n2097;
  assign n2391 = n2390 ^ n2094;
  assign n2392 = ~n2095 & n2391;
  assign n2393 = n2392 ^ n2094;
  assign n2394 = n2393 ^ n2089;
  assign n2395 = ~n2090 & n2394;
  assign n2396 = n2395 ^ n2087;
  assign n2397 = n2396 ^ n2084;
  assign n2398 = ~n2085 & ~n2397;
  assign n2399 = n2398 ^ n2084;
  assign n2400 = n2399 ^ n2077;
  assign n2401 = ~n2078 & ~n2400;
  assign n2402 = n2401 ^ n2074;
  assign n2403 = n2402 ^ n2070;
  assign n2404 = ~n2071 & n2403;
  assign n2405 = n2404 ^ n2068;
  assign n2406 = n2405 ^ n2065;
  assign n2407 = ~n2066 & ~n2406;
  assign n2408 = n2407 ^ n2065;
  assign n2409 = n2408 ^ n2060;
  assign n2410 = ~n2061 & ~n2409;
  assign n2411 = n2410 ^ n2060;
  assign n2412 = n2411 ^ n2050;
  assign n2413 = ~n2054 & ~n2412;
  assign n2414 = n2413 ^ n2053;
  assign n2415 = n2414 ^ n2046;
  assign n2416 = ~n2047 & ~n2415;
  assign n2417 = n2416 ^ n2044;
  assign n2418 = n2417 ^ n2041;
  assign n2419 = ~n2042 & ~n2418;
  assign n2420 = n2419 ^ n2041;
  assign n2421 = n2420 ^ n2036;
  assign n2422 = ~n2037 & ~n2421;
  assign n2423 = n2422 ^ n2033;
  assign n2424 = n2423 ^ n2029;
  assign n2425 = ~n2030 & n2424;
  assign n2426 = n2425 ^ n2029;
  assign n2427 = n2426 ^ n2022;
  assign n2428 = ~n2023 & ~n2427;
  assign n2429 = n2428 ^ n2022;
  assign n2430 = n2429 ^ n2013;
  assign n2431 = ~n2017 & ~n2430;
  assign n2432 = n2431 ^ n2013;
  assign n2433 = n2432 ^ n2010;
  assign n2434 = ~n2011 & ~n2433;
  assign n2435 = n2434 ^ n2008;
  assign n2436 = n2435 ^ n2004;
  assign n2437 = ~n2005 & ~n2436;
  assign n2438 = n2437 ^ n2002;
  assign n2439 = n2438 ^ n1999;
  assign n2440 = ~n2000 & n2439;
  assign n2441 = n2440 ^ n1999;
  assign n2442 = n2441 ^ n1994;
  assign n2443 = ~n1995 & ~n2442;
  assign n2444 = n2443 ^ n1994;
  assign n2445 = n2444 ^ n1987;
  assign n2446 = ~n1990 & n2445;
  assign n2447 = n2446 ^ n1989;
  assign n2448 = n2447 ^ n1984;
  assign n2449 = ~n1985 & ~n2448;
  assign n2450 = n2449 ^ n1982;
  assign n2451 = n2450 ^ n1979;
  assign n2452 = ~n1980 & n2451;
  assign n2453 = n2452 ^ n1979;
  assign n2454 = n2453 ^ n1974;
  assign n2455 = ~n1975 & n2454;
  assign n2456 = n2455 ^ n1974;
  assign n2457 = n2456 ^ n1966;
  assign n2458 = ~n1970 & n2457;
  assign n2459 = n2458 ^ n1966;
  assign n2460 = n2459 ^ n1962;
  assign n2461 = ~n1963 & ~n2460;
  assign n2462 = n2461 ^ n1962;
  assign n2463 = n2462 ^ n1952;
  assign n2464 = ~n1956 & ~n2463;
  assign n2465 = n2464 ^ n1952;
  assign n2466 = n2465 ^ n1949;
  assign n2467 = ~n1950 & ~n2466;
  assign n2468 = n2467 ^ n1949;
  assign n2469 = n2468 ^ n1940;
  assign n2470 = ~n1944 & n2469;
  assign n2471 = n2470 ^ n1940;
  assign n2472 = n2471 ^ n1937;
  assign n2473 = ~n1938 & n2472;
  assign n2474 = n2473 ^ n1937;
  assign n2475 = n2474 ^ n1929;
  assign n2476 = ~n1932 & n2475;
  assign n2477 = n2476 ^ n1929;
  assign n2478 = n2477 ^ n1926;
  assign n2479 = ~n1927 & ~n2478;
  assign n2480 = n2479 ^ n1924;
  assign n2481 = n2480 ^ n1921;
  assign n2482 = ~n1922 & n2481;
  assign n2483 = n2482 ^ n1918;
  assign n2484 = n2483 ^ n1915;
  assign n2485 = ~n1916 & n2484;
  assign n2486 = n2485 ^ n1915;
  assign n2487 = n2486 ^ n1908;
  assign n2488 = ~n1909 & ~n2487;
  assign n2489 = n2488 ^ n1908;
  assign n2490 = n2489 ^ n1901;
  assign n2491 = ~n1904 & ~n2490;
  assign n2492 = n2491 ^ n1903;
  assign n2493 = n2492 ^ n1898;
  assign n2494 = ~n1899 & n2493;
  assign n2495 = n2494 ^ n1895;
  assign n2496 = n2495 ^ n1891;
  assign n2497 = ~n1892 & ~n2496;
  assign n2498 = n2497 ^ n1891;
  assign n2499 = n2498 ^ n1885;
  assign n2500 = ~n1886 & ~n2499;
  assign n2501 = n2500 ^ n1885;
  assign n2502 = n2501 ^ n1879;
  assign n2503 = ~n1880 & n2502;
  assign n2504 = n2503 ^ n1879;
  assign n2505 = n2504 ^ n1870;
  assign n2506 = ~n1874 & ~n2505;
  assign n2507 = n2506 ^ n1870;
  assign n2508 = n2507 ^ n1867;
  assign n2509 = ~n1868 & ~n2508;
  assign n2510 = n2509 ^ n1867;
  assign n2511 = n2510 ^ n1859;
  assign n2512 = ~n1862 & ~n2511;
  assign n2513 = n2512 ^ n1861;
  assign n2514 = n2513 ^ n1855;
  assign n2515 = ~n1856 & n2514;
  assign n2516 = n2515 ^ n1852;
  assign n2517 = n2516 ^ n1847;
  assign n2518 = ~n1850 & ~n2517;
  assign n2519 = n2518 ^ n1847;
  assign n2520 = n2519 ^ n1843;
  assign n2521 = ~n1844 & n2520;
  assign n2522 = n2521 ^ n1841;
  assign n2523 = n2522 ^ n1837;
  assign n2524 = ~n1838 & n2523;
  assign n2525 = n2524 ^ n1835;
  assign n2526 = n2525 ^ n1830;
  assign n2527 = ~n1833 & ~n2526;
  assign n2528 = n2527 ^ n1830;
  assign n2529 = n2528 ^ n1825;
  assign n2530 = ~n1828 & ~n2529;
  assign n2531 = n2530 ^ n1825;
  assign n2532 = n2531 ^ n1822;
  assign n2533 = ~n1823 & n2532;
  assign n2534 = n2533 ^ n1822;
  assign n2535 = n2534 ^ n1815;
  assign n2536 = ~n1818 & n2535;
  assign n2537 = n2536 ^ n1815;
  assign n2538 = n2537 ^ n1810;
  assign n2539 = ~n1813 & n2538;
  assign n2540 = n2539 ^ n1810;
  assign n2541 = n2540 ^ n1805;
  assign n2542 = ~n1808 & n2541;
  assign n2543 = n2542 ^ n1805;
  assign n2544 = n2543 ^ n1802;
  assign n2545 = ~n1803 & ~n2544;
  assign n2546 = n2545 ^ n1802;
  assign n2547 = n2546 ^ n1795;
  assign n2548 = ~n1798 & n2547;
  assign n2549 = n2548 ^ n1795;
  assign n2550 = n2549 ^ n1792;
  assign n2551 = ~n1793 & n2550;
  assign n2552 = n2551 ^ n1792;
  assign n2553 = n2552 ^ n1785;
  assign n2554 = ~n1788 & ~n2553;
  assign n2555 = n2554 ^ n1785;
  assign n2556 = n2555 ^ n1780;
  assign n2557 = ~n1783 & ~n2556;
  assign n2558 = n2557 ^ n1782;
  assign n2559 = n2558 ^ n1777;
  assign n2560 = ~n1778 & n2559;
  assign n2561 = n2560 ^ n1775;
  assign n2562 = n2561 ^ n1770;
  assign n2563 = ~n1773 & n2562;
  assign n2564 = n2563 ^ n1770;
  assign n2565 = n2564 ^ n1765;
  assign n2566 = ~n1768 & n2565;
  assign n2567 = n2566 ^ n1765;
  assign n2568 = n2567 ^ n1760;
  assign n2569 = ~n1763 & ~n2568;
  assign n2570 = n2569 ^ n1762;
  assign n2571 = n2570 ^ n1757;
  assign n2572 = ~n1758 & n2571;
  assign n2573 = n2572 ^ n1755;
  assign n2574 = n2573 ^ n1750;
  assign n2575 = ~n1753 & ~n2574;
  assign n2576 = n2575 ^ n1750;
  assign n2577 = n2576 ^ n1745;
  assign n2578 = ~n1748 & n2577;
  assign n2579 = n2578 ^ n1745;
  assign n2580 = n2579 ^ n1742;
  assign n2581 = ~n1743 & ~n2580;
  assign n2582 = n2581 ^ n1740;
  assign n2583 = n2582 ^ n1737;
  assign n2584 = ~n1738 & n2583;
  assign n2585 = n2584 ^ n1735;
  assign n2586 = n2585 ^ n1730;
  assign n2587 = ~n1733 & ~n2586;
  assign n2588 = n2587 ^ n1730;
  assign n2589 = n2588 ^ n1725;
  assign n2590 = ~n1728 & n2589;
  assign n2591 = n2590 ^ n1727;
  assign n2592 = n2591 ^ n1722;
  assign n2593 = ~n1723 & ~n2592;
  assign n2594 = n2593 ^ n1720;
  assign n2595 = n2594 ^ n1715;
  assign n2596 = ~n1718 & ~n2595;
  assign n2597 = n2596 ^ n1715;
  assign n2598 = n2597 ^ n1712;
  assign n2599 = ~n1713 & n2598;
  assign n2600 = n2599 ^ n1710;
  assign n2601 = n2600 ^ n1707;
  assign n2602 = ~n1708 & n2601;
  assign n2603 = n2602 ^ n1705;
  assign n2604 = n2603 ^ n1702;
  assign n2605 = ~n1703 & n2604;
  assign n2606 = n2605 ^ n1702;
  assign n2607 = n2606 ^ n1697;
  assign n2608 = ~n1698 & ~n2607;
  assign n2609 = n2608 ^ n1695;
  assign n2610 = n2609 ^ n1692;
  assign n2611 = ~n1693 & n2610;
  assign n2612 = n2611 ^ n1690;
  assign n2613 = n2612 ^ n1685;
  assign n2614 = ~n1688 & ~n2613;
  assign n2615 = n2614 ^ n1685;
  assign n2616 = n2615 ^ n1680;
  assign n2617 = ~n1683 & n2616;
  assign n2618 = n2617 ^ n1680;
  assign n2619 = n2618 ^ n1677;
  assign n2620 = ~n1678 & ~n2619;
  assign n2621 = n2620 ^ n1677;
  assign n2622 = n2621 ^ n1670;
  assign n2623 = ~n1673 & ~n2622;
  assign n2624 = n2623 ^ n1670;
  assign n2625 = n2624 ^ n1667;
  assign n2626 = ~n1668 & n2625;
  assign n2627 = n2626 ^ n1667;
  assign n2628 = n2627 ^ n1660;
  assign n2629 = ~n1663 & ~n2628;
  assign n2630 = n2629 ^ n1660;
  assign n2631 = n2630 ^ n1657;
  assign n2632 = ~n1658 & n2631;
  assign n2633 = n2632 ^ n1657;
  assign n2634 = n2633 ^ n1652;
  assign n2635 = ~n1653 & ~n2634;
  assign n2636 = n2635 ^ n1650;
  assign n2637 = n2636 ^ n1647;
  assign n2638 = ~n1648 & n2637;
  assign n2639 = n2638 ^ n1645;
  assign n2640 = n2639 ^ n1642;
  assign n2641 = ~n1643 & n2640;
  assign n2642 = n2641 ^ n1642;
  assign n2643 = n2642 ^ n1635;
  assign n2644 = ~n1638 & ~n2643;
  assign n2645 = n2644 ^ n1637;
  assign n2646 = n2645 ^ n1632;
  assign n2647 = ~n1633 & ~n2646;
  assign n2648 = n2647 ^ n1630;
  assign n2649 = n2648 ^ n1624;
  assign n2650 = ~n1628 & n2649;
  assign n2651 = n2650 ^ n1624;
  assign n2652 = n2651 ^ n1617;
  assign n2653 = ~n1621 & n2652;
  assign n2654 = n2653 ^ n1617;
  assign n2655 = n2654 ^ n1613;
  assign n2656 = ~n1614 & ~n2655;
  assign n2657 = n2656 ^ n1613;
  assign n2658 = n2657 ^ n1062;
  assign n2659 = ~n1609 & ~n2658;
  assign n2661 = n2660 ^ n2659;
  assign n2662 = ~n515 & n2661;
  assign n2663 = n2662 ^ n513;
  assign n2664 = n2281 ^ n2278;
  assign n2665 = ~n2663 & n2664;
  assign n2666 = n2665 ^ n2278;
  assign n2667 = n2275 & ~n2663;
  assign n2668 = n2667 ^ n2272;
  assign n2669 = n2270 & ~n2663;
  assign n2670 = n2669 ^ n2267;
  assign n2671 = n2265 & ~n2663;
  assign n2672 = n2671 ^ n2264;
  assign n2673 = n2260 & n2663;
  assign n2674 = n2673 ^ n2257;
  assign n2675 = n2255 & n2663;
  assign n2676 = n2675 ^ n2252;
  assign n2677 = n2250 & ~n2663;
  assign n2678 = n2677 ^ n2247;
  assign n2679 = n2245 & n2663;
  assign n2680 = n2679 ^ n2242;
  assign n2681 = n2240 & ~n2663;
  assign n2682 = n2681 ^ n2237;
  assign n2683 = n2235 & ~n2663;
  assign n2684 = n2683 ^ n2232;
  assign n2685 = n2230 & n2663;
  assign n2686 = n2685 ^ n2229;
  assign n2687 = n2225 & n2663;
  assign n2688 = n2687 ^ n2222;
  assign n2689 = n2220 & n2663;
  assign n2690 = n2689 ^ n2219;
  assign n2691 = n2215 & ~n2663;
  assign n2692 = n2691 ^ n2212;
  assign n2693 = n2210 & ~n2663;
  assign n2694 = n2693 ^ n2209;
  assign n2695 = n2205 & n2663;
  assign n2696 = n2695 ^ n2202;
  assign n2697 = n2200 & ~n2663;
  assign n2698 = n2697 ^ n2197;
  assign n2699 = n2195 & n2663;
  assign n2700 = n2699 ^ n2192;
  assign n2701 = n2190 & n2663;
  assign n2702 = n2701 ^ n2187;
  assign n2703 = n2185 & ~n2663;
  assign n2704 = n2703 ^ n2182;
  assign n2705 = n2180 & n2663;
  assign n2706 = n2705 ^ n2177;
  assign n2707 = n2175 & ~n2663;
  assign n2708 = n2707 ^ n2172;
  assign n2709 = n2170 & ~n2663;
  assign n2710 = n2709 ^ n2167;
  assign n2711 = n2165 & ~n2663;
  assign n2712 = n2711 ^ n2164;
  assign n2713 = n2160 & n2663;
  assign n2714 = n2713 ^ n2157;
  assign n2715 = n2155 & n2663;
  assign n2716 = n2715 ^ n2152;
  assign n2717 = n2150 & n2663;
  assign n2718 = n2717 ^ n2147;
  assign n2719 = n2145 & ~n2663;
  assign n2720 = n2719 ^ n2142;
  assign n2721 = n2140 & n2663;
  assign n2722 = n2721 ^ n2137;
  assign n2723 = n2135 & n2663;
  assign n2724 = n2723 ^ n2132;
  assign n2725 = n2130 & ~n2663;
  assign n2726 = n2725 ^ n2127;
  assign n2727 = n2125 & n2663;
  assign n2728 = n2727 ^ n2122;
  assign n2729 = n2120 & n2663;
  assign n2730 = n2729 ^ n2117;
  assign n2731 = n2115 & n2663;
  assign n2732 = n2731 ^ n2112;
  assign n2733 = n2110 & ~n2663;
  assign n2734 = n2733 ^ n2107;
  assign n2735 = n2105 & n2663;
  assign n2736 = n2735 ^ n2104;
  assign n2737 = n2100 & n2663;
  assign n2738 = n2737 ^ n2097;
  assign n2739 = n2095 & ~n2663;
  assign n2740 = n2739 ^ n2092;
  assign n2741 = n2090 & n2663;
  assign n2742 = n2741 ^ n2087;
  assign n2743 = n2085 & n2663;
  assign n2744 = n2743 ^ n2081;
  assign n2745 = n2078 & n2663;
  assign n2746 = n2745 ^ n2074;
  assign n2747 = n2071 & n2663;
  assign n2748 = n2747 ^ n2068;
  assign n2749 = n2066 & n2663;
  assign n2750 = n2749 ^ n2063;
  assign n2751 = n2061 & ~n2663;
  assign n2752 = n2751 ^ n2057;
  assign n2753 = n2054 & ~n2663;
  assign n2754 = n2753 ^ n2053;
  assign n2755 = n2047 & n2663;
  assign n2756 = n2755 ^ n2044;
  assign n2757 = n2042 & n2663;
  assign n2758 = n2757 ^ n2039;
  assign n2759 = n2037 & n2663;
  assign n2760 = n2759 ^ n2033;
  assign n2761 = n2030 & ~n2663;
  assign n2762 = n2761 ^ n2026;
  assign n2763 = n2023 & n2663;
  assign n2764 = n2763 ^ n2019;
  assign n2765 = n2017 & ~n2663;
  assign n2766 = n2765 ^ n2016;
  assign n2767 = n2011 & ~n2663;
  assign n2768 = n2767 ^ n2008;
  assign n2769 = n2005 & n2663;
  assign n2770 = n2769 ^ n2002;
  assign n2771 = n2000 & ~n2663;
  assign n2772 = n2771 ^ n1997;
  assign n2773 = n1995 & n2663;
  assign n2774 = n2773 ^ n1992;
  assign n2775 = n1990 & ~n2663;
  assign n2776 = n2775 ^ n1989;
  assign n2777 = n1985 & n2663;
  assign n2778 = n2777 ^ n1982;
  assign n2779 = n1980 & ~n2663;
  assign n2780 = n2779 ^ n1977;
  assign n2781 = n1975 & ~n2663;
  assign n2782 = n2781 ^ n1972;
  assign n2783 = n1970 & ~n2663;
  assign n2784 = n2783 ^ n1969;
  assign n2785 = n1963 & n2663;
  assign n2786 = n2785 ^ n1959;
  assign n2787 = n1956 & ~n2663;
  assign n2788 = n2787 ^ n1955;
  assign n2789 = n1950 & n2663;
  assign n2790 = n2789 ^ n1946;
  assign n2791 = n1944 & n2663;
  assign n2792 = n2791 ^ n1943;
  assign n2793 = n1938 & n2663;
  assign n2794 = n2793 ^ n1934;
  assign n2795 = n1932 & n2663;
  assign n2796 = n2795 ^ n1931;
  assign n2797 = n1927 & n2663;
  assign n2798 = n2797 ^ n1924;
  assign n2799 = n1922 & n2663;
  assign n2800 = n2799 ^ n1918;
  assign n2801 = n1916 & ~n2663;
  assign n2802 = n2801 ^ n1912;
  assign n2803 = n1909 & n2663;
  assign n2804 = n2803 ^ n1906;
  assign n2805 = n1904 & n2663;
  assign n2806 = n2805 ^ n1903;
  assign n2807 = n1899 & n2663;
  assign n2808 = n2807 ^ n1895;
  assign n2809 = n1892 & n2663;
  assign n2810 = n2809 ^ n1889;
  assign n2811 = n1886 & ~n2663;
  assign n2812 = n2811 ^ n1882;
  assign n2813 = n1880 & n2663;
  assign n2814 = n2813 ^ n1879;
  assign n2815 = n1874 & ~n2663;
  assign n2816 = n2815 ^ n1870;
  assign n2817 = n1868 & n2663;
  assign n2818 = n2817 ^ n1867;
  assign n2819 = n1862 & ~n2663;
  assign n2820 = n2819 ^ n1861;
  assign n2821 = n1856 & ~n2663;
  assign n2822 = n2821 ^ n1852;
  assign n2823 = n1850 & n2663;
  assign n2824 = n2823 ^ n1847;
  assign n2825 = n1844 & n2663;
  assign n2826 = n2825 ^ n1841;
  assign n2827 = n1838 & n2663;
  assign n2828 = n2827 ^ n1835;
  assign n2829 = n1833 & ~n2663;
  assign n2830 = n2829 ^ n1830;
  assign n2831 = n1828 & n2663;
  assign n2832 = n2831 ^ n1825;
  assign n2833 = n1823 & n2663;
  assign n2834 = n2833 ^ n1822;
  assign n2835 = n1818 & n2663;
  assign n2836 = n2835 ^ n1815;
  assign n2837 = n1813 & ~n2663;
  assign n2838 = n2837 ^ n1812;
  assign n2839 = n1808 & n2663;
  assign n2840 = n2839 ^ n1805;
  assign n2841 = n1803 & ~n2663;
  assign n2842 = n2841 ^ n1802;
  assign n2843 = n1798 & ~n2663;
  assign n2844 = n2843 ^ n1795;
  assign n2845 = n1793 & ~n2663;
  assign n2846 = n2845 ^ n1792;
  assign n2847 = n1788 & n2663;
  assign n2848 = n2847 ^ n1785;
  assign n2849 = n1783 & ~n2663;
  assign n2850 = n2849 ^ n1782;
  assign n2851 = n1778 & ~n2663;
  assign n2852 = n2851 ^ n1775;
  assign n2853 = n1773 & ~n2663;
  assign n2854 = n2853 ^ n1770;
  assign n2855 = n1768 & ~n2663;
  assign n2856 = n2855 ^ n1765;
  assign n2857 = n1763 & n2663;
  assign n2858 = n2857 ^ n1762;
  assign n2859 = n1758 & n2663;
  assign n2860 = n2859 ^ n1755;
  assign n2861 = n1753 & ~n2663;
  assign n2862 = n2861 ^ n1750;
  assign n2863 = n1748 & ~n2663;
  assign n2864 = n2863 ^ n1745;
  assign n2865 = n1743 & n2663;
  assign n2866 = n2865 ^ n1740;
  assign n2867 = n1738 & n2663;
  assign n2868 = n2867 ^ n1735;
  assign n2869 = n1733 & ~n2663;
  assign n2870 = n2869 ^ n1730;
  assign n2871 = n1728 & ~n2663;
  assign n2872 = n2871 ^ n1727;
  assign n2873 = n1723 & n2663;
  assign n2874 = n2873 ^ n1720;
  assign n2875 = n1718 & ~n2663;
  assign n2876 = n2875 ^ n1715;
  assign n2877 = n1713 & ~n2663;
  assign n2878 = n2877 ^ n1710;
  assign n2879 = n1708 & ~n2663;
  assign n2880 = n2879 ^ n1705;
  assign n2881 = n1703 & n2663;
  assign n2882 = n2881 ^ n1700;
  assign n2883 = n1698 & n2663;
  assign n2884 = n2883 ^ n1695;
  assign n2885 = n1693 & n2663;
  assign n2886 = n2885 ^ n1690;
  assign n2887 = n1688 & ~n2663;
  assign n2888 = n2887 ^ n1685;
  assign n2889 = n1683 & ~n2663;
  assign n2890 = n2889 ^ n1680;
  assign n2891 = n1678 & n2663;
  assign n2892 = n2891 ^ n1677;
  assign n2893 = n1673 & ~n2663;
  assign n2894 = n2893 ^ n1670;
  assign n2895 = n1668 & ~n2663;
  assign n2896 = n2895 ^ n1667;
  assign n2897 = n1663 & n2663;
  assign n2898 = n2897 ^ n1660;
  assign n2899 = n1658 & n2663;
  assign n2900 = n2899 ^ n1657;
  assign n2901 = n1653 & ~n2663;
  assign n2902 = n2901 ^ n1650;
  assign n2903 = n1648 & ~n2663;
  assign n2904 = n2903 ^ n1645;
  assign n2905 = n1643 & n2663;
  assign n2906 = n2905 ^ n1640;
  assign n2907 = n1638 & n2663;
  assign n2908 = n2907 ^ n1637;
  assign n2909 = n1633 & ~n2663;
  assign n2910 = n2909 ^ n1630;
  assign n2911 = n1628 & ~n2663;
  assign n2912 = n2911 ^ n1624;
  assign n2913 = n1621 & ~n2663;
  assign n2914 = n2913 ^ n1617;
  assign n2915 = n1614 & n2663;
  assign n2916 = n2915 ^ n1613;
  assign n2917 = n1609 & ~n2663;
  assign n2918 = n2917 ^ n1608;
  assign n2919 = n513 & n514;
  assign n2920 = n1606 ^ n1060;
  assign n2921 = ~n2663 & n2920;
  assign n2922 = n2921 ^ n1606;
  assign y0 = n2666;
  assign y1 = n2668;
  assign y2 = n2670;
  assign y3 = n2672;
  assign y4 = n2674;
  assign y5 = n2676;
  assign y6 = n2678;
  assign y7 = n2680;
  assign y8 = n2682;
  assign y9 = n2684;
  assign y10 = n2686;
  assign y11 = n2688;
  assign y12 = n2690;
  assign y13 = n2692;
  assign y14 = n2694;
  assign y15 = n2696;
  assign y16 = n2698;
  assign y17 = n2700;
  assign y18 = n2702;
  assign y19 = n2704;
  assign y20 = n2706;
  assign y21 = n2708;
  assign y22 = n2710;
  assign y23 = n2712;
  assign y24 = n2714;
  assign y25 = n2716;
  assign y26 = n2718;
  assign y27 = n2720;
  assign y28 = n2722;
  assign y29 = n2724;
  assign y30 = n2726;
  assign y31 = n2728;
  assign y32 = n2730;
  assign y33 = n2732;
  assign y34 = n2734;
  assign y35 = n2736;
  assign y36 = n2738;
  assign y37 = n2740;
  assign y38 = n2742;
  assign y39 = n2744;
  assign y40 = n2746;
  assign y41 = n2748;
  assign y42 = n2750;
  assign y43 = n2752;
  assign y44 = n2754;
  assign y45 = n2756;
  assign y46 = n2758;
  assign y47 = n2760;
  assign y48 = n2762;
  assign y49 = n2764;
  assign y50 = n2766;
  assign y51 = n2768;
  assign y52 = n2770;
  assign y53 = n2772;
  assign y54 = n2774;
  assign y55 = n2776;
  assign y56 = n2778;
  assign y57 = n2780;
  assign y58 = n2782;
  assign y59 = n2784;
  assign y60 = n2786;
  assign y61 = n2788;
  assign y62 = n2790;
  assign y63 = n2792;
  assign y64 = n2794;
  assign y65 = n2796;
  assign y66 = n2798;
  assign y67 = n2800;
  assign y68 = n2802;
  assign y69 = n2804;
  assign y70 = n2806;
  assign y71 = n2808;
  assign y72 = n2810;
  assign y73 = n2812;
  assign y74 = n2814;
  assign y75 = n2816;
  assign y76 = n2818;
  assign y77 = n2820;
  assign y78 = n2822;
  assign y79 = n2824;
  assign y80 = n2826;
  assign y81 = n2828;
  assign y82 = n2830;
  assign y83 = n2832;
  assign y84 = n2834;
  assign y85 = n2836;
  assign y86 = n2838;
  assign y87 = n2840;
  assign y88 = n2842;
  assign y89 = n2844;
  assign y90 = n2846;
  assign y91 = n2848;
  assign y92 = n2850;
  assign y93 = n2852;
  assign y94 = n2854;
  assign y95 = n2856;
  assign y96 = n2858;
  assign y97 = n2860;
  assign y98 = n2862;
  assign y99 = n2864;
  assign y100 = n2866;
  assign y101 = n2868;
  assign y102 = n2870;
  assign y103 = n2872;
  assign y104 = n2874;
  assign y105 = n2876;
  assign y106 = n2878;
  assign y107 = n2880;
  assign y108 = n2882;
  assign y109 = n2884;
  assign y110 = n2886;
  assign y111 = n2888;
  assign y112 = n2890;
  assign y113 = n2892;
  assign y114 = n2894;
  assign y115 = n2896;
  assign y116 = n2898;
  assign y117 = n2900;
  assign y118 = n2902;
  assign y119 = n2904;
  assign y120 = n2906;
  assign y121 = n2908;
  assign y122 = n2910;
  assign y123 = n2912;
  assign y124 = n2914;
  assign y125 = n2916;
  assign y126 = n2918;
  assign y127 = n2919;
  assign y128 = n2922;
  assign y129 = n2663;
endmodule